***********************PLL-final*****************************

.param L=0.15
.param W=0.42

