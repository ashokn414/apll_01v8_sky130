magic
tech sky130A
timestamp 1605505535
<< nwell >>
rect -20 -190 1500 90
<< nmos >>
rect 100 -411 115 -369
rect 270 -411 285 -369
rect 315 -411 330 -369
rect 480 -411 495 -369
rect 525 -411 540 -369
rect 690 -411 705 -369
rect 735 -411 750 -369
rect 900 -411 915 -369
rect 945 -411 960 -369
rect 1110 -411 1125 -369
rect 1155 -411 1170 -369
rect 1320 -411 1335 -369
<< pmos >>
rect 100 -134 115 -50
rect 270 -134 285 -50
rect 315 -134 330 -50
rect 480 -134 495 -50
rect 525 -134 540 -50
rect 690 -134 705 -50
rect 735 -134 750 -50
rect 900 -134 915 -50
rect 945 -134 960 -50
rect 1110 -134 1125 -50
rect 1155 -134 1170 -50
rect 1320 -134 1335 -50
<< ndiff >>
rect 40 -377 100 -369
rect 40 -401 48 -377
rect 72 -401 100 -377
rect 40 -411 100 -401
rect 115 -377 170 -369
rect 115 -401 138 -377
rect 162 -401 170 -377
rect 115 -411 170 -401
rect 210 -377 270 -369
rect 210 -401 218 -377
rect 242 -401 270 -377
rect 210 -411 270 -401
rect 285 -411 315 -369
rect 330 -377 380 -369
rect 330 -401 348 -377
rect 372 -401 380 -377
rect 330 -411 380 -401
rect 420 -377 480 -369
rect 420 -401 428 -377
rect 452 -401 480 -377
rect 420 -411 480 -401
rect 495 -411 525 -369
rect 540 -377 590 -369
rect 540 -401 558 -377
rect 582 -401 590 -377
rect 540 -411 590 -401
rect 630 -377 690 -369
rect 630 -401 638 -377
rect 662 -401 690 -377
rect 630 -411 690 -401
rect 705 -411 735 -369
rect 750 -377 800 -369
rect 750 -401 768 -377
rect 792 -401 800 -377
rect 750 -411 800 -401
rect 840 -377 900 -369
rect 840 -401 848 -377
rect 872 -401 900 -377
rect 840 -411 900 -401
rect 915 -411 945 -369
rect 960 -377 1010 -369
rect 960 -401 978 -377
rect 1002 -401 1010 -377
rect 960 -411 1010 -401
rect 1050 -377 1110 -369
rect 1050 -401 1058 -377
rect 1082 -401 1110 -377
rect 1050 -411 1110 -401
rect 1125 -411 1155 -369
rect 1170 -377 1220 -369
rect 1170 -401 1188 -377
rect 1212 -401 1220 -377
rect 1170 -411 1220 -401
rect 1260 -377 1320 -369
rect 1260 -401 1268 -377
rect 1292 -401 1320 -377
rect 1260 -411 1320 -401
rect 1335 -377 1390 -369
rect 1335 -401 1358 -377
rect 1382 -401 1390 -377
rect 1335 -411 1390 -401
<< pdiff >>
rect 40 -76 100 -50
rect 40 -106 47 -76
rect 77 -106 100 -76
rect 40 -134 100 -106
rect 115 -76 170 -50
rect 115 -106 133 -76
rect 163 -106 170 -76
rect 115 -134 170 -106
rect 210 -76 270 -50
rect 210 -106 217 -76
rect 247 -106 270 -76
rect 210 -134 270 -106
rect 285 -134 315 -50
rect 330 -76 380 -50
rect 330 -106 343 -76
rect 373 -106 380 -76
rect 330 -134 380 -106
rect 420 -76 480 -50
rect 420 -106 427 -76
rect 457 -106 480 -76
rect 420 -134 480 -106
rect 495 -134 525 -50
rect 540 -76 590 -50
rect 540 -106 553 -76
rect 583 -106 590 -76
rect 540 -134 590 -106
rect 630 -76 690 -50
rect 630 -106 637 -76
rect 667 -106 690 -76
rect 630 -134 690 -106
rect 705 -134 735 -50
rect 750 -76 800 -50
rect 750 -106 763 -76
rect 793 -106 800 -76
rect 750 -134 800 -106
rect 840 -76 900 -50
rect 840 -106 847 -76
rect 877 -106 900 -76
rect 840 -134 900 -106
rect 915 -134 945 -50
rect 960 -76 1010 -50
rect 960 -106 973 -76
rect 1003 -106 1010 -76
rect 960 -134 1010 -106
rect 1050 -76 1110 -50
rect 1050 -106 1057 -76
rect 1087 -106 1110 -76
rect 1050 -134 1110 -106
rect 1125 -134 1155 -50
rect 1170 -76 1220 -50
rect 1170 -106 1183 -76
rect 1213 -106 1220 -76
rect 1170 -134 1220 -106
rect 1260 -76 1320 -50
rect 1260 -106 1267 -76
rect 1297 -106 1320 -76
rect 1260 -134 1320 -106
rect 1335 -76 1390 -50
rect 1335 -106 1353 -76
rect 1383 -106 1390 -76
rect 1335 -134 1390 -106
<< ndiffc >>
rect 48 -401 72 -377
rect 138 -401 162 -377
rect 218 -401 242 -377
rect 348 -401 372 -377
rect 428 -401 452 -377
rect 558 -401 582 -377
rect 638 -401 662 -377
rect 768 -401 792 -377
rect 848 -401 872 -377
rect 978 -401 1002 -377
rect 1058 -401 1082 -377
rect 1188 -401 1212 -377
rect 1268 -401 1292 -377
rect 1358 -401 1382 -377
<< pdiffc >>
rect 47 -106 77 -76
rect 133 -106 163 -76
rect 217 -106 247 -76
rect 343 -106 373 -76
rect 427 -106 457 -76
rect 553 -106 583 -76
rect 637 -106 667 -76
rect 763 -106 793 -76
rect 847 -106 877 -76
rect 973 -106 1003 -76
rect 1057 -106 1087 -76
rect 1183 -106 1213 -76
rect 1267 -106 1297 -76
rect 1353 -106 1383 -76
<< psubdiff >>
rect 0 -489 1460 -479
rect 0 -529 20 -489
rect 60 -529 111 -489
rect 151 -529 200 -489
rect 240 -529 291 -489
rect 331 -529 414 -489
rect 455 -529 516 -489
rect 556 -529 620 -489
rect 660 -529 718 -489
rect 758 -529 834 -489
rect 875 -529 921 -489
rect 961 -529 1040 -489
rect 1080 -529 1146 -489
rect 1186 -529 1251 -489
rect 1292 -529 1326 -489
rect 1366 -529 1400 -489
rect 1440 -529 1460 -489
rect 0 -539 1460 -529
<< nsubdiff >>
rect 0 60 1480 70
rect 0 20 20 60
rect 60 20 140 60
rect 180 20 260 60
rect 300 20 380 60
rect 420 20 500 60
rect 540 20 620 60
rect 660 20 740 60
rect 780 20 860 60
rect 900 20 1000 60
rect 1040 20 1120 60
rect 1160 20 1240 60
rect 1280 20 1360 60
rect 1400 20 1480 60
rect 0 10 1480 20
<< psubdiffcont >>
rect 20 -529 60 -489
rect 111 -529 151 -489
rect 200 -529 240 -489
rect 291 -529 331 -489
rect 414 -529 455 -489
rect 516 -529 556 -489
rect 620 -529 660 -489
rect 718 -529 758 -489
rect 834 -529 875 -489
rect 921 -529 961 -489
rect 1040 -529 1080 -489
rect 1146 -529 1186 -489
rect 1251 -529 1292 -489
rect 1326 -529 1366 -489
rect 1400 -529 1440 -489
<< nsubdiffcont >>
rect 20 20 60 60
rect 140 20 180 60
rect 260 20 300 60
rect 380 20 420 60
rect 500 20 540 60
rect 620 20 660 60
rect 740 20 780 60
rect 860 20 900 60
rect 1000 20 1040 60
rect 1120 20 1160 60
rect 1240 20 1280 60
rect 1360 20 1400 60
<< poly >>
rect 100 -50 115 -30
rect 270 -50 285 -30
rect 315 -50 330 -30
rect 480 -50 495 -30
rect 525 -50 540 -30
rect 690 -50 705 -30
rect 735 -50 750 -30
rect 900 -50 915 -30
rect 945 -50 960 -30
rect 1110 -50 1125 -30
rect 1155 -50 1170 -30
rect 1320 -50 1335 -30
rect 100 -160 115 -134
rect 270 -160 285 -134
rect 100 -170 140 -160
rect 100 -190 110 -170
rect 130 -190 140 -170
rect 100 -200 140 -190
rect 245 -170 285 -160
rect 245 -190 255 -170
rect 275 -190 285 -170
rect 245 -200 285 -190
rect 315 -227 330 -134
rect 480 -160 495 -134
rect 455 -170 495 -160
rect 455 -190 465 -170
rect 485 -190 495 -170
rect 455 -200 495 -190
rect 280 -237 330 -227
rect 525 -230 540 -134
rect 690 -160 705 -134
rect 665 -170 705 -160
rect 665 -190 675 -170
rect 695 -190 705 -170
rect 665 -200 705 -190
rect 735 -230 750 -134
rect 900 -160 915 -134
rect 875 -170 915 -160
rect 875 -190 885 -170
rect 905 -190 915 -170
rect 875 -200 915 -190
rect 945 -230 960 -134
rect 1110 -160 1125 -134
rect 1085 -170 1125 -160
rect 1085 -190 1095 -170
rect 1115 -190 1125 -170
rect 1085 -200 1125 -190
rect 1155 -230 1170 -134
rect 1320 -230 1335 -134
rect 280 -268 291 -237
rect 320 -268 330 -237
rect 280 -277 330 -268
rect 500 -240 540 -230
rect 500 -260 510 -240
rect 530 -260 540 -240
rect 500 -270 540 -260
rect 710 -240 750 -230
rect 710 -260 720 -240
rect 740 -260 750 -240
rect 710 -270 750 -260
rect 920 -240 960 -230
rect 920 -260 930 -240
rect 950 -260 960 -240
rect 920 -270 960 -260
rect 1130 -240 1170 -230
rect 1130 -260 1140 -240
rect 1160 -260 1170 -240
rect 1130 -270 1170 -260
rect 80 -309 120 -299
rect 80 -329 90 -309
rect 110 -329 120 -309
rect 80 -339 120 -329
rect 250 -309 290 -299
rect 250 -329 260 -309
rect 280 -329 290 -309
rect 250 -339 290 -329
rect 100 -369 115 -339
rect 270 -369 285 -339
rect 315 -369 330 -277
rect 460 -309 500 -299
rect 460 -329 470 -309
rect 490 -329 500 -309
rect 460 -339 500 -329
rect 480 -369 495 -339
rect 525 -369 540 -270
rect 670 -309 710 -299
rect 670 -329 680 -309
rect 700 -329 710 -309
rect 670 -339 710 -329
rect 690 -369 705 -339
rect 735 -369 750 -270
rect 880 -309 920 -299
rect 880 -329 890 -309
rect 910 -329 920 -309
rect 880 -339 920 -329
rect 900 -369 915 -339
rect 945 -369 960 -270
rect 1090 -309 1130 -299
rect 1090 -329 1100 -309
rect 1120 -329 1130 -309
rect 1090 -339 1130 -329
rect 1110 -369 1125 -339
rect 1155 -369 1170 -270
rect 1290 -242 1335 -230
rect 1290 -263 1302 -242
rect 1324 -263 1335 -242
rect 1290 -274 1335 -263
rect 1320 -369 1335 -274
rect 100 -429 115 -411
rect 270 -429 285 -411
rect 315 -429 330 -411
rect 480 -429 495 -411
rect 525 -429 540 -411
rect 690 -429 705 -411
rect 735 -429 750 -411
rect 900 -429 915 -411
rect 945 -429 960 -411
rect 1110 -429 1125 -411
rect 1155 -429 1170 -411
rect 1320 -429 1335 -411
<< polycont >>
rect 110 -190 130 -170
rect 255 -190 275 -170
rect 465 -190 485 -170
rect 675 -190 695 -170
rect 885 -190 905 -170
rect 1095 -190 1115 -170
rect 291 -268 320 -237
rect 510 -260 530 -240
rect 720 -260 740 -240
rect 930 -260 950 -240
rect 1140 -260 1160 -240
rect 90 -329 110 -309
rect 260 -329 280 -309
rect 470 -329 490 -309
rect 680 -329 700 -309
rect 890 -329 910 -309
rect 1100 -329 1120 -309
rect 1302 -263 1324 -242
<< locali >>
rect 0 60 1480 80
rect 0 20 20 60
rect 60 20 140 60
rect 180 20 260 60
rect 300 20 380 60
rect 420 20 500 60
rect 540 20 620 60
rect 660 20 740 60
rect 780 20 860 60
rect 900 20 1000 60
rect 1040 20 1120 60
rect 1160 20 1240 60
rect 1280 20 1360 60
rect 1400 20 1480 60
rect 0 0 1480 20
rect 40 -50 70 0
rect 210 -50 240 0
rect 420 -50 450 0
rect 630 -50 660 0
rect 840 -50 870 0
rect 1050 -50 1080 0
rect 1260 -50 1290 0
rect 40 -76 80 -50
rect 40 -106 47 -76
rect 77 -106 80 -76
rect 40 -134 80 -106
rect 130 -76 170 -50
rect 130 -106 133 -76
rect 163 -106 170 -76
rect 130 -134 170 -106
rect 210 -76 250 -50
rect 210 -106 217 -76
rect 247 -106 250 -76
rect 210 -134 250 -106
rect 340 -76 380 -50
rect 340 -106 343 -76
rect 373 -106 380 -76
rect 340 -134 380 -106
rect 420 -76 460 -50
rect 420 -106 427 -76
rect 457 -106 460 -76
rect 420 -134 460 -106
rect 550 -76 590 -50
rect 550 -106 553 -76
rect 583 -106 590 -76
rect 550 -134 590 -106
rect 630 -76 670 -50
rect 630 -106 637 -76
rect 667 -106 670 -76
rect 630 -134 670 -106
rect 760 -76 800 -50
rect 760 -106 763 -76
rect 793 -106 800 -76
rect 760 -134 800 -106
rect 840 -76 880 -50
rect 840 -106 847 -76
rect 877 -106 880 -76
rect 840 -134 880 -106
rect 970 -76 1010 -50
rect 970 -106 973 -76
rect 1003 -106 1010 -76
rect 970 -134 1010 -106
rect 1050 -76 1090 -50
rect 1050 -106 1057 -76
rect 1087 -106 1090 -76
rect 1050 -134 1090 -106
rect 1180 -76 1220 -50
rect 1180 -106 1183 -76
rect 1213 -106 1220 -76
rect 1180 -134 1220 -106
rect 1260 -76 1300 -50
rect 1260 -106 1267 -76
rect 1297 -106 1300 -76
rect 1260 -134 1300 -106
rect 1350 -76 1390 -50
rect 1350 -106 1353 -76
rect 1383 -106 1390 -76
rect 1350 -134 1390 -106
rect 140 -160 170 -134
rect 100 -170 170 -160
rect 100 -190 110 -170
rect 130 -190 170 -170
rect 100 -200 170 -190
rect 245 -170 285 -160
rect 245 -190 255 -170
rect 275 -190 285 -170
rect 245 -200 285 -190
rect 80 -309 120 -299
rect 40 -329 90 -309
rect 110 -329 120 -309
rect 40 -339 120 -329
rect 140 -369 170 -200
rect 280 -237 330 -227
rect 280 -268 291 -237
rect 320 -268 330 -237
rect 280 -277 330 -268
rect 350 -240 380 -134
rect 455 -170 495 -160
rect 455 -190 465 -170
rect 485 -190 495 -170
rect 455 -200 495 -190
rect 500 -240 540 -230
rect 350 -260 510 -240
rect 530 -260 540 -240
rect 350 -270 540 -260
rect 560 -240 590 -134
rect 665 -170 705 -160
rect 665 -190 675 -170
rect 695 -190 705 -170
rect 665 -200 705 -190
rect 710 -240 750 -230
rect 560 -260 720 -240
rect 740 -260 750 -240
rect 560 -270 750 -260
rect 770 -240 800 -134
rect 875 -170 915 -160
rect 875 -190 885 -170
rect 905 -190 915 -170
rect 875 -200 915 -190
rect 920 -240 960 -230
rect 770 -260 930 -240
rect 950 -260 960 -240
rect 770 -270 960 -260
rect 980 -240 1010 -134
rect 1085 -170 1125 -160
rect 1085 -190 1095 -170
rect 1115 -190 1125 -170
rect 1085 -200 1125 -190
rect 1190 -230 1220 -134
rect 1130 -240 1170 -230
rect 980 -260 1140 -240
rect 1160 -260 1170 -240
rect 980 -270 1170 -260
rect 1190 -240 1240 -230
rect 1290 -240 1335 -230
rect 1360 -240 1390 -134
rect 1190 -270 1200 -240
rect 1230 -242 1335 -240
rect 1230 -263 1302 -242
rect 1324 -263 1335 -242
rect 1230 -270 1335 -263
rect 1359 -270 1450 -240
rect 250 -309 290 -299
rect 250 -329 260 -309
rect 280 -329 290 -309
rect 250 -339 290 -329
rect 350 -369 380 -270
rect 460 -309 500 -299
rect 460 -329 470 -309
rect 490 -329 500 -309
rect 460 -339 500 -329
rect 560 -369 590 -270
rect 670 -309 710 -299
rect 670 -329 680 -309
rect 700 -329 710 -309
rect 670 -339 710 -329
rect 770 -369 800 -270
rect 880 -309 920 -299
rect 880 -329 890 -309
rect 910 -329 920 -309
rect 880 -339 920 -329
rect 980 -369 1010 -270
rect 1190 -280 1240 -270
rect 1290 -274 1335 -270
rect 1090 -309 1130 -299
rect 1090 -329 1100 -309
rect 1120 -329 1130 -309
rect 1090 -339 1130 -329
rect 1190 -369 1220 -280
rect 1360 -369 1390 -270
rect 40 -377 80 -369
rect 40 -401 48 -377
rect 72 -401 80 -377
rect 40 -411 80 -401
rect 130 -377 170 -369
rect 130 -401 138 -377
rect 162 -401 170 -377
rect 130 -411 170 -401
rect 210 -377 250 -369
rect 210 -401 218 -377
rect 242 -401 250 -377
rect 210 -411 250 -401
rect 340 -377 380 -369
rect 340 -401 348 -377
rect 372 -401 380 -377
rect 340 -411 380 -401
rect 420 -377 460 -369
rect 420 -401 428 -377
rect 452 -401 460 -377
rect 420 -411 460 -401
rect 550 -377 590 -369
rect 550 -401 558 -377
rect 582 -401 590 -377
rect 550 -411 590 -401
rect 630 -377 670 -369
rect 630 -401 638 -377
rect 662 -401 670 -377
rect 630 -411 670 -401
rect 760 -377 800 -369
rect 760 -401 768 -377
rect 792 -401 800 -377
rect 760 -411 800 -401
rect 840 -377 880 -369
rect 840 -401 848 -377
rect 872 -401 880 -377
rect 840 -411 880 -401
rect 970 -377 1010 -369
rect 970 -401 978 -377
rect 1002 -401 1010 -377
rect 970 -411 1010 -401
rect 1050 -377 1090 -369
rect 1050 -401 1058 -377
rect 1082 -401 1090 -377
rect 1050 -411 1090 -401
rect 1180 -377 1220 -369
rect 1180 -401 1188 -377
rect 1212 -401 1220 -377
rect 1180 -411 1220 -401
rect 1260 -377 1300 -369
rect 1260 -401 1268 -377
rect 1292 -401 1300 -377
rect 1260 -411 1300 -401
rect 1350 -377 1390 -369
rect 1350 -401 1358 -377
rect 1382 -401 1390 -377
rect 1350 -411 1390 -401
rect 40 -469 70 -411
rect 210 -469 240 -411
rect 420 -469 450 -411
rect 630 -469 660 -411
rect 840 -469 870 -411
rect 1050 -469 1080 -411
rect 1260 -469 1290 -411
rect 0 -489 1460 -469
rect 0 -529 20 -489
rect 60 -529 111 -489
rect 151 -529 200 -489
rect 240 -529 291 -489
rect 331 -529 414 -489
rect 455 -529 516 -489
rect 556 -529 620 -489
rect 660 -529 718 -489
rect 758 -529 834 -489
rect 875 -529 921 -489
rect 961 -529 1040 -489
rect 1080 -529 1146 -489
rect 1186 -529 1251 -489
rect 1292 -529 1326 -489
rect 1366 -529 1400 -489
rect 1440 -529 1460 -489
rect 0 -549 1460 -529
<< viali >>
rect 110 -190 130 -170
rect 255 -190 275 -170
rect 90 -329 110 -309
rect 291 -268 320 -237
rect 465 -190 485 -170
rect 675 -190 695 -170
rect 885 -190 905 -170
rect 1095 -190 1115 -170
rect 1200 -270 1230 -240
rect 260 -329 280 -309
rect 470 -329 490 -309
rect 680 -329 700 -309
rect 890 -329 910 -309
rect 1100 -329 1120 -309
<< metal1 >>
rect 100 -170 140 -160
rect 245 -170 285 -160
rect 455 -170 495 -160
rect 665 -170 705 -160
rect 875 -170 915 -160
rect 1085 -170 1125 -160
rect 100 -190 110 -170
rect 130 -190 255 -170
rect 275 -190 465 -170
rect 485 -190 675 -170
rect 695 -190 885 -170
rect 905 -190 1095 -170
rect 1115 -190 1125 -170
rect 100 -200 1125 -190
rect 280 -237 330 -227
rect 280 -268 291 -237
rect 320 -268 330 -237
rect 280 -277 330 -268
rect 1190 -240 1240 -230
rect 1190 -270 1200 -240
rect 1230 -270 1240 -240
rect 1190 -280 1240 -270
rect 80 -309 120 -299
rect 250 -309 290 -299
rect 460 -309 500 -299
rect 670 -309 710 -299
rect 880 -309 920 -299
rect 1090 -309 1130 -299
rect 80 -329 90 -309
rect 110 -329 260 -309
rect 280 -329 470 -309
rect 490 -329 680 -309
rect 700 -329 890 -309
rect 910 -329 1100 -309
rect 1120 -329 1130 -309
rect 80 -339 1130 -329
<< via1 >>
rect 291 -268 320 -237
rect 1200 -270 1230 -240
<< metal2 >>
rect 280 -237 330 -227
rect 280 -268 291 -237
rect 320 -268 330 -237
rect 280 -277 330 -268
rect 1190 -240 1240 -230
rect 1190 -270 1200 -240
rect 1230 -270 1240 -240
rect 1190 -280 1240 -270
<< via2 >>
rect 291 -268 320 -237
rect 1200 -270 1230 -240
<< metal3 >>
rect 280 -230 330 -227
rect 280 -237 1240 -230
rect 280 -268 291 -237
rect 320 -240 1240 -237
rect 320 -268 1200 -240
rect 280 -270 1200 -268
rect 1230 -270 1240 -240
rect 280 -277 330 -270
rect 1190 -280 1240 -270
<< labels >>
rlabel locali 688 36 720 52 1 vdd
rlabel locali 706 -524 738 -508 1 gnd!
rlabel locali 48 -330 71 -320 1 vin
rlabel locali 1419 -260 1442 -250 1 vout
<< end >>
