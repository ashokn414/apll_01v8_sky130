magic
tech sky130A
timestamp 1605604810
<< nwell >>
rect -130 -290 1245 30
rect -130 -410 1246 -290
rect -130 -1871 1263 -1491
<< nmos >>
rect 40 438 55 480
rect 200 396 215 480
rect 280 396 295 480
rect 440 438 455 480
rect 600 438 615 480
rect 760 354 775 480
rect 840 354 855 480
rect 925 354 940 480
rect 1120 438 1135 480
rect 340 -916 355 -832
rect 425 -916 440 -832
rect 600 -916 615 -832
rect 685 -916 700 -832
rect 860 -916 875 -748
rect 940 -916 955 -748
rect 1020 -916 1035 -748
rect 1100 -916 1115 -748
rect 340 -1180 355 -1096
rect 425 -1180 440 -1096
rect 600 -1180 615 -1096
rect 685 -1180 700 -1096
rect 37 -2311 52 -2269
rect 197 -2311 212 -2227
rect 277 -2311 292 -2227
rect 437 -2311 452 -2269
rect 597 -2311 612 -2269
rect 790 -2311 805 -2185
rect 870 -2311 885 -2185
rect 955 -2311 970 -2185
rect 1150 -2311 1165 -2269
<< pmos >>
rect 40 -80 55 4
rect 200 -80 215 4
rect 280 -80 295 4
rect 440 -80 455 4
rect 600 -80 615 4
rect 760 -80 775 4
rect 840 -80 855 4
rect 925 -80 940 4
rect 1120 -80 1135 4
rect 340 -384 355 -300
rect 425 -384 440 -300
rect 600 -384 615 -300
rect 685 -384 700 -300
rect 860 -384 875 -300
rect 940 -384 955 -300
rect 1020 -384 1035 -300
rect 1100 -384 1115 -300
rect 340 -1601 355 -1517
rect 425 -1601 440 -1517
rect 600 -1601 615 -1517
rect 685 -1601 700 -1517
rect 37 -1845 52 -1761
rect 197 -1845 212 -1761
rect 277 -1845 292 -1761
rect 437 -1845 452 -1761
rect 597 -1845 612 -1761
rect 790 -1845 805 -1761
rect 870 -1845 885 -1761
rect 955 -1845 970 -1761
rect 1150 -1845 1165 -1761
<< ndiff >>
rect -10 472 40 480
rect -10 448 -2 472
rect 22 448 40 472
rect -10 438 40 448
rect 55 472 110 480
rect 55 448 78 472
rect 102 448 110 472
rect 55 438 110 448
rect 150 473 200 480
rect 150 405 158 473
rect 182 405 200 473
rect 150 396 200 405
rect 215 396 280 480
rect 295 472 345 480
rect 295 404 313 472
rect 337 404 345 472
rect 390 472 440 480
rect 390 448 398 472
rect 422 448 440 472
rect 390 438 440 448
rect 455 472 510 480
rect 455 448 478 472
rect 502 448 510 472
rect 455 438 510 448
rect 550 472 600 480
rect 550 448 558 472
rect 582 448 600 472
rect 550 438 600 448
rect 615 472 670 480
rect 615 448 638 472
rect 662 448 670 472
rect 615 438 670 448
rect 710 452 760 480
rect 295 396 345 404
rect 710 384 718 452
rect 742 384 760 452
rect 710 354 760 384
rect 775 354 840 480
rect 855 354 925 480
rect 940 445 990 480
rect 940 377 958 445
rect 982 377 990 445
rect 1070 472 1120 480
rect 1070 448 1078 472
rect 1102 448 1120 472
rect 1070 438 1120 448
rect 1135 472 1190 480
rect 1135 448 1158 472
rect 1182 448 1190 472
rect 1135 438 1190 448
rect 940 354 990 377
rect 810 -780 860 -748
rect 290 -840 340 -832
rect 290 -908 298 -840
rect 322 -908 340 -840
rect 290 -916 340 -908
rect 355 -916 425 -832
rect 440 -840 490 -832
rect 440 -908 458 -840
rect 482 -908 490 -840
rect 440 -916 490 -908
rect 550 -840 600 -832
rect 550 -908 558 -840
rect 582 -908 600 -840
rect 550 -916 600 -908
rect 615 -916 685 -832
rect 700 -840 750 -832
rect 700 -908 718 -840
rect 742 -908 750 -840
rect 700 -916 750 -908
rect 810 -899 818 -780
rect 841 -899 860 -780
rect 810 -916 860 -899
rect 875 -916 940 -748
rect 955 -916 1020 -748
rect 1035 -916 1100 -748
rect 1115 -776 1171 -748
rect 1115 -897 1137 -776
rect 1163 -897 1171 -776
rect 1115 -916 1171 -897
rect 1129 -917 1171 -916
rect 450 -1096 492 -1094
rect 290 -1104 340 -1096
rect 290 -1172 298 -1104
rect 322 -1172 340 -1104
rect 290 -1180 340 -1172
rect 355 -1180 425 -1096
rect 440 -1104 492 -1096
rect 440 -1172 458 -1104
rect 484 -1172 492 -1104
rect 440 -1180 492 -1172
rect 550 -1104 600 -1096
rect 550 -1172 558 -1104
rect 582 -1172 600 -1104
rect 550 -1180 600 -1172
rect 615 -1180 685 -1096
rect 700 -1104 750 -1096
rect 700 -1172 718 -1104
rect 742 -1172 750 -1104
rect 700 -1180 750 -1172
rect 147 -2235 197 -2227
rect -13 -2279 37 -2269
rect -13 -2303 -5 -2279
rect 19 -2303 37 -2279
rect -13 -2311 37 -2303
rect 52 -2279 107 -2269
rect 52 -2303 75 -2279
rect 99 -2303 107 -2279
rect 52 -2311 107 -2303
rect 147 -2303 155 -2235
rect 179 -2303 197 -2235
rect 147 -2311 197 -2303
rect 212 -2311 277 -2227
rect 292 -2235 342 -2227
rect 292 -2303 311 -2235
rect 335 -2303 342 -2235
rect 740 -2221 790 -2185
rect 292 -2311 342 -2303
rect 387 -2279 437 -2269
rect 387 -2303 395 -2279
rect 419 -2303 437 -2279
rect 387 -2311 437 -2303
rect 452 -2279 507 -2269
rect 452 -2303 475 -2279
rect 499 -2303 507 -2279
rect 452 -2311 507 -2303
rect 547 -2279 597 -2269
rect 547 -2303 555 -2279
rect 579 -2303 597 -2279
rect 547 -2311 597 -2303
rect 612 -2279 667 -2269
rect 612 -2303 635 -2279
rect 659 -2303 667 -2279
rect 612 -2311 667 -2303
rect 740 -2289 748 -2221
rect 772 -2289 790 -2221
rect 740 -2311 790 -2289
rect 805 -2311 870 -2185
rect 885 -2311 955 -2185
rect 970 -2212 1020 -2185
rect 970 -2280 988 -2212
rect 1012 -2280 1020 -2212
rect 970 -2311 1020 -2280
rect 1100 -2279 1150 -2269
rect 1100 -2303 1108 -2279
rect 1132 -2303 1150 -2279
rect 1100 -2311 1150 -2303
rect 1165 -2279 1220 -2269
rect 1165 -2303 1188 -2279
rect 1212 -2303 1220 -2279
rect 1165 -2311 1220 -2303
<< pdiff >>
rect -10 -20 40 4
rect -10 -60 -4 -20
rect 26 -60 40 -20
rect -10 -80 40 -60
rect 55 -20 110 4
rect 55 -60 73 -20
rect 103 -60 110 -20
rect 55 -80 110 -60
rect 150 -20 200 4
rect 150 -60 156 -20
rect 186 -60 200 -20
rect 150 -80 200 -60
rect 215 -20 280 4
rect 215 -60 232 -20
rect 262 -60 280 -20
rect 215 -80 280 -60
rect 295 -20 345 4
rect 295 -60 310 -20
rect 340 -60 345 -20
rect 295 -80 345 -60
rect 390 -20 440 4
rect 390 -60 396 -20
rect 426 -60 440 -20
rect 390 -80 440 -60
rect 455 -20 510 4
rect 455 -60 473 -20
rect 503 -60 510 -20
rect 455 -80 510 -60
rect 550 -20 600 4
rect 550 -60 556 -20
rect 586 -60 600 -20
rect 550 -80 600 -60
rect 615 -20 670 4
rect 615 -60 633 -20
rect 663 -60 670 -20
rect 615 -80 670 -60
rect 710 -20 760 4
rect 710 -60 716 -20
rect 746 -60 760 -20
rect 710 -80 760 -60
rect 775 -20 840 4
rect 775 -60 794 -20
rect 824 -60 840 -20
rect 775 -80 840 -60
rect 855 -20 925 4
rect 855 -60 876 -20
rect 906 -60 925 -20
rect 855 -80 925 -60
rect 940 -20 990 4
rect 940 -60 955 -20
rect 985 -60 990 -20
rect 940 -80 990 -60
rect 1070 -20 1120 4
rect 1070 -60 1076 -20
rect 1106 -60 1120 -20
rect 1070 -80 1120 -60
rect 1135 -20 1190 4
rect 1135 -60 1153 -20
rect 1183 -60 1190 -20
rect 1135 -80 1190 -60
rect 290 -320 340 -300
rect 290 -360 296 -320
rect 326 -360 340 -320
rect 290 -384 340 -360
rect 355 -320 425 -300
rect 355 -360 375 -320
rect 405 -360 425 -320
rect 355 -384 425 -360
rect 440 -320 490 -300
rect 440 -360 453 -320
rect 483 -360 490 -320
rect 440 -384 490 -360
rect 550 -320 600 -300
rect 550 -360 556 -320
rect 586 -360 600 -320
rect 550 -384 600 -360
rect 615 -320 685 -300
rect 615 -360 635 -320
rect 665 -360 685 -320
rect 615 -384 685 -360
rect 700 -320 750 -300
rect 700 -360 713 -320
rect 743 -360 750 -320
rect 700 -384 750 -360
rect 810 -319 860 -300
rect 810 -359 816 -319
rect 846 -359 860 -319
rect 810 -384 860 -359
rect 875 -320 940 -300
rect 875 -360 895 -320
rect 925 -360 940 -320
rect 875 -384 940 -360
rect 955 -319 1020 -300
rect 955 -359 976 -319
rect 1006 -359 1020 -319
rect 955 -384 1020 -359
rect 1035 -319 1100 -300
rect 1035 -359 1056 -319
rect 1086 -359 1100 -319
rect 1035 -384 1100 -359
rect 1115 -319 1170 -300
rect 1115 -359 1136 -319
rect 1166 -359 1170 -319
rect 1115 -384 1170 -359
rect 290 -1541 340 -1517
rect 290 -1581 296 -1541
rect 326 -1581 340 -1541
rect 290 -1601 340 -1581
rect 355 -1541 425 -1517
rect 355 -1581 375 -1541
rect 405 -1581 425 -1541
rect 355 -1601 425 -1581
rect 440 -1541 490 -1517
rect 440 -1581 453 -1541
rect 483 -1581 490 -1541
rect 440 -1601 490 -1581
rect 550 -1541 600 -1517
rect 550 -1581 556 -1541
rect 586 -1581 600 -1541
rect 550 -1601 600 -1581
rect 615 -1541 685 -1517
rect 615 -1581 635 -1541
rect 665 -1581 685 -1541
rect 615 -1601 685 -1581
rect 700 -1541 750 -1517
rect 700 -1581 713 -1541
rect 743 -1581 750 -1541
rect 700 -1601 750 -1581
rect -13 -1781 37 -1761
rect -13 -1821 -7 -1781
rect 23 -1821 37 -1781
rect -13 -1845 37 -1821
rect 52 -1781 107 -1761
rect 52 -1821 70 -1781
rect 100 -1821 107 -1781
rect 52 -1845 107 -1821
rect 147 -1781 197 -1761
rect 147 -1821 153 -1781
rect 183 -1821 197 -1781
rect 147 -1845 197 -1821
rect 212 -1781 277 -1761
rect 212 -1821 229 -1781
rect 259 -1821 277 -1781
rect 212 -1845 277 -1821
rect 292 -1781 342 -1761
rect 292 -1821 307 -1781
rect 337 -1821 342 -1781
rect 292 -1845 342 -1821
rect 387 -1781 437 -1761
rect 387 -1821 393 -1781
rect 423 -1821 437 -1781
rect 387 -1845 437 -1821
rect 452 -1781 507 -1761
rect 452 -1821 470 -1781
rect 500 -1821 507 -1781
rect 452 -1845 507 -1821
rect 547 -1781 597 -1761
rect 547 -1821 553 -1781
rect 583 -1821 597 -1781
rect 547 -1845 597 -1821
rect 612 -1781 667 -1761
rect 612 -1821 630 -1781
rect 660 -1821 667 -1781
rect 612 -1845 667 -1821
rect 740 -1781 790 -1761
rect 740 -1821 745 -1781
rect 776 -1821 790 -1781
rect 740 -1845 790 -1821
rect 805 -1781 870 -1761
rect 805 -1821 824 -1781
rect 854 -1821 870 -1781
rect 805 -1845 870 -1821
rect 885 -1781 955 -1761
rect 885 -1821 906 -1781
rect 936 -1821 955 -1781
rect 885 -1845 955 -1821
rect 970 -1781 1020 -1761
rect 970 -1821 985 -1781
rect 1015 -1821 1020 -1781
rect 970 -1845 1020 -1821
rect 1100 -1781 1150 -1761
rect 1100 -1821 1106 -1781
rect 1136 -1821 1150 -1781
rect 1100 -1845 1150 -1821
rect 1165 -1781 1220 -1761
rect 1165 -1821 1183 -1781
rect 1213 -1821 1220 -1781
rect 1165 -1845 1220 -1821
<< ndiffc >>
rect -2 448 22 472
rect 78 448 102 472
rect 158 405 182 473
rect 313 404 337 472
rect 398 448 422 472
rect 478 448 502 472
rect 558 448 582 472
rect 638 448 662 472
rect 718 384 742 452
rect 958 377 982 445
rect 1078 448 1102 472
rect 1158 448 1182 472
rect 298 -908 322 -840
rect 458 -908 482 -840
rect 558 -908 582 -840
rect 718 -908 742 -840
rect 818 -899 841 -780
rect 1137 -897 1163 -776
rect 298 -1172 322 -1104
rect 458 -1172 484 -1104
rect 558 -1172 582 -1104
rect 718 -1172 742 -1104
rect -5 -2303 19 -2279
rect 75 -2303 99 -2279
rect 155 -2303 179 -2235
rect 311 -2303 335 -2235
rect 395 -2303 419 -2279
rect 475 -2303 499 -2279
rect 555 -2303 579 -2279
rect 635 -2303 659 -2279
rect 748 -2289 772 -2221
rect 988 -2280 1012 -2212
rect 1108 -2303 1132 -2279
rect 1188 -2303 1212 -2279
<< pdiffc >>
rect -4 -60 26 -20
rect 73 -60 103 -20
rect 156 -60 186 -20
rect 232 -60 262 -20
rect 310 -60 340 -20
rect 396 -60 426 -20
rect 473 -60 503 -20
rect 556 -60 586 -20
rect 633 -60 663 -20
rect 716 -60 746 -20
rect 794 -60 824 -20
rect 876 -60 906 -20
rect 955 -60 985 -20
rect 1076 -60 1106 -20
rect 1153 -60 1183 -20
rect 296 -360 326 -320
rect 375 -360 405 -320
rect 453 -360 483 -320
rect 556 -360 586 -320
rect 635 -360 665 -320
rect 713 -360 743 -320
rect 816 -359 846 -319
rect 895 -360 925 -320
rect 976 -359 1006 -319
rect 1056 -359 1086 -319
rect 1136 -359 1166 -319
rect 296 -1581 326 -1541
rect 375 -1581 405 -1541
rect 453 -1581 483 -1541
rect 556 -1581 586 -1541
rect 635 -1581 665 -1541
rect 713 -1581 743 -1541
rect -7 -1821 23 -1781
rect 70 -1821 100 -1781
rect 153 -1821 183 -1781
rect 229 -1821 259 -1781
rect 307 -1821 337 -1781
rect 393 -1821 423 -1781
rect 470 -1821 500 -1781
rect 553 -1821 583 -1781
rect 630 -1821 660 -1781
rect 745 -1821 776 -1781
rect 824 -1821 854 -1781
rect 906 -1821 936 -1781
rect 985 -1821 1015 -1781
rect 1106 -1821 1136 -1781
rect 1183 -1821 1213 -1781
<< psubdiff >>
rect -60 590 1380 600
rect -60 550 -40 590
rect 0 550 40 590
rect 80 550 120 590
rect 160 550 200 590
rect 240 550 280 590
rect 320 550 360 590
rect 400 550 440 590
rect 480 550 520 590
rect 560 550 600 590
rect 640 550 680 590
rect 720 550 760 590
rect 800 550 840 590
rect 880 550 920 590
rect 960 550 1000 590
rect 1040 550 1080 590
rect 1120 550 1160 590
rect 1200 550 1240 590
rect 1280 550 1320 590
rect 1360 550 1380 590
rect -60 540 1380 550
rect 1320 530 1380 540
rect 1320 490 1330 530
rect 1370 490 1380 530
rect 1320 450 1380 490
rect 1320 310 1330 450
rect 1370 310 1380 450
rect 1320 270 1380 310
rect 1320 230 1330 270
rect 1370 230 1380 270
rect 1320 190 1380 230
rect 1320 150 1330 190
rect 1370 150 1380 190
rect 1320 110 1380 150
rect 1320 70 1330 110
rect 1370 70 1380 110
rect 1320 30 1380 70
rect 1320 -10 1330 30
rect 1370 -10 1380 30
rect 1320 -50 1380 -10
rect 1320 -90 1330 -50
rect 1370 -90 1380 -50
rect 1320 -130 1380 -90
rect 1320 -170 1330 -130
rect 1370 -170 1380 -130
rect 1320 -210 1380 -170
rect 1320 -250 1330 -210
rect 1370 -250 1380 -210
rect 1320 -290 1380 -250
rect 1320 -330 1330 -290
rect 1370 -330 1380 -290
rect 1320 -370 1380 -330
rect 1320 -410 1330 -370
rect 1370 -410 1380 -370
rect 1320 -450 1380 -410
rect 1320 -490 1330 -450
rect 1370 -490 1380 -450
rect 1320 -530 1380 -490
rect 1320 -570 1330 -530
rect 1370 -570 1380 -530
rect 1320 -610 1380 -570
rect 1320 -650 1330 -610
rect 1370 -650 1380 -610
rect 1320 -690 1380 -650
rect 1320 -886 1330 -690
rect 1370 -886 1380 -690
rect 1320 -926 1380 -886
rect 1320 -966 1330 -926
rect 1370 -966 1380 -926
rect 1320 -976 1380 -966
rect 290 -986 1380 -976
rect 290 -1026 310 -986
rect 350 -1026 390 -986
rect 430 -1026 830 -986
rect 870 -1026 910 -986
rect 950 -1026 990 -986
rect 1030 -1026 1070 -986
rect 1110 -1026 1270 -986
rect 1310 -1006 1380 -986
rect 1310 -1026 1330 -1006
rect 290 -1036 1330 -1026
rect 1320 -1046 1330 -1036
rect 1370 -1046 1380 -1006
rect 1320 -1086 1380 -1046
rect 1320 -1126 1330 -1086
rect 1370 -1126 1380 -1086
rect 1320 -1211 1380 -1126
rect 1320 -1251 1330 -1211
rect 1370 -1251 1380 -1211
rect 1320 -1291 1380 -1251
rect 1320 -1331 1330 -1291
rect 1370 -1331 1380 -1291
rect 1320 -1371 1380 -1331
rect 1320 -1411 1330 -1371
rect 1370 -1411 1380 -1371
rect 1320 -1451 1380 -1411
rect 1320 -1491 1330 -1451
rect 1370 -1491 1380 -1451
rect 1320 -1531 1380 -1491
rect 1320 -1571 1330 -1531
rect 1370 -1571 1380 -1531
rect 1320 -1611 1380 -1571
rect 1320 -1651 1330 -1611
rect 1370 -1651 1380 -1611
rect 1320 -1691 1380 -1651
rect 1320 -1731 1330 -1691
rect 1370 -1731 1380 -1691
rect 1320 -1771 1380 -1731
rect 1320 -1811 1330 -1771
rect 1370 -1811 1380 -1771
rect 1320 -1851 1380 -1811
rect 1320 -1891 1330 -1851
rect 1370 -1891 1380 -1851
rect 1320 -1931 1380 -1891
rect 1320 -1971 1330 -1931
rect 1370 -1971 1380 -1931
rect 1320 -2011 1380 -1971
rect 1320 -2051 1330 -2011
rect 1370 -2051 1380 -2011
rect 1320 -2091 1380 -2051
rect 1320 -2131 1330 -2091
rect 1370 -2131 1380 -2091
rect 1320 -2261 1380 -2131
rect 1320 -2301 1330 -2261
rect 1370 -2301 1380 -2261
rect 1320 -2371 1380 -2301
rect -60 -2381 1330 -2371
rect -60 -2421 -40 -2381
rect 0 -2421 40 -2381
rect 80 -2421 120 -2381
rect 160 -2421 200 -2381
rect 240 -2421 280 -2381
rect 320 -2421 360 -2381
rect 400 -2421 440 -2381
rect 480 -2421 520 -2381
rect 560 -2421 600 -2381
rect 640 -2421 680 -2381
rect 720 -2421 760 -2381
rect 800 -2421 840 -2381
rect 880 -2421 920 -2381
rect 960 -2421 1000 -2381
rect 1040 -2421 1080 -2381
rect 1120 -2421 1160 -2381
rect 1200 -2421 1240 -2381
rect 1280 -2411 1330 -2381
rect 1370 -2411 1380 -2371
rect 1280 -2421 1380 -2411
rect -60 -2431 1380 -2421
<< nsubdiff >>
rect -90 -140 1220 -130
rect -90 -180 -50 -140
rect -10 -180 20 -140
rect 60 -180 90 -140
rect 130 -180 160 -140
rect 200 -180 310 -140
rect 350 -180 740 -140
rect 780 -180 800 -140
rect 840 -180 870 -140
rect 910 -180 940 -140
rect 980 -180 1100 -140
rect 1140 -180 1160 -140
rect 1200 -180 1220 -140
rect -90 -190 1220 -180
rect -90 -1661 1230 -1651
rect -90 -1701 -70 -1661
rect -30 -1701 0 -1661
rect 40 -1701 70 -1661
rect 110 -1701 140 -1661
rect 180 -1701 300 -1661
rect 340 -1701 750 -1661
rect 790 -1701 820 -1661
rect 860 -1701 890 -1661
rect 930 -1701 960 -1661
rect 1000 -1701 1100 -1661
rect 1140 -1701 1170 -1661
rect 1210 -1701 1230 -1661
rect -90 -1711 1230 -1701
<< psubdiffcont >>
rect -40 550 0 590
rect 40 550 80 590
rect 120 550 160 590
rect 200 550 240 590
rect 280 550 320 590
rect 360 550 400 590
rect 440 550 480 590
rect 520 550 560 590
rect 600 550 640 590
rect 680 550 720 590
rect 760 550 800 590
rect 840 550 880 590
rect 920 550 960 590
rect 1000 550 1040 590
rect 1080 550 1120 590
rect 1160 550 1200 590
rect 1240 550 1280 590
rect 1320 550 1360 590
rect 1330 490 1370 530
rect 1330 310 1370 450
rect 1330 230 1370 270
rect 1330 150 1370 190
rect 1330 70 1370 110
rect 1330 -10 1370 30
rect 1330 -90 1370 -50
rect 1330 -170 1370 -130
rect 1330 -250 1370 -210
rect 1330 -330 1370 -290
rect 1330 -410 1370 -370
rect 1330 -490 1370 -450
rect 1330 -570 1370 -530
rect 1330 -650 1370 -610
rect 1330 -886 1370 -690
rect 1330 -966 1370 -926
rect 310 -1026 350 -986
rect 390 -1026 430 -986
rect 830 -1026 870 -986
rect 910 -1026 950 -986
rect 990 -1026 1030 -986
rect 1070 -1026 1110 -986
rect 1270 -1026 1310 -986
rect 1330 -1046 1370 -1006
rect 1330 -1126 1370 -1086
rect 1330 -1251 1370 -1211
rect 1330 -1331 1370 -1291
rect 1330 -1411 1370 -1371
rect 1330 -1491 1370 -1451
rect 1330 -1571 1370 -1531
rect 1330 -1651 1370 -1611
rect 1330 -1731 1370 -1691
rect 1330 -1811 1370 -1771
rect 1330 -1891 1370 -1851
rect 1330 -1971 1370 -1931
rect 1330 -2051 1370 -2011
rect 1330 -2131 1370 -2091
rect 1330 -2301 1370 -2261
rect -40 -2421 0 -2381
rect 40 -2421 80 -2381
rect 120 -2421 160 -2381
rect 200 -2421 240 -2381
rect 280 -2421 320 -2381
rect 360 -2421 400 -2381
rect 440 -2421 480 -2381
rect 520 -2421 560 -2381
rect 600 -2421 640 -2381
rect 680 -2421 720 -2381
rect 760 -2421 800 -2381
rect 840 -2421 880 -2381
rect 920 -2421 960 -2381
rect 1000 -2421 1040 -2381
rect 1080 -2421 1120 -2381
rect 1160 -2421 1200 -2381
rect 1240 -2421 1280 -2381
rect 1330 -2411 1370 -2371
<< nsubdiffcont >>
rect -50 -180 -10 -140
rect 20 -180 60 -140
rect 90 -180 130 -140
rect 160 -180 200 -140
rect 310 -180 350 -140
rect 740 -180 780 -140
rect 800 -180 840 -140
rect 870 -180 910 -140
rect 940 -180 980 -140
rect 1100 -180 1140 -140
rect 1160 -180 1200 -140
rect -70 -1701 -30 -1661
rect 0 -1701 40 -1661
rect 70 -1701 110 -1661
rect 140 -1701 180 -1661
rect 300 -1701 340 -1661
rect 750 -1701 790 -1661
rect 820 -1701 860 -1661
rect 890 -1701 930 -1661
rect 960 -1701 1000 -1661
rect 1100 -1701 1140 -1661
rect 1170 -1701 1210 -1661
<< poly >>
rect 40 480 55 500
rect 200 480 215 500
rect 280 480 295 500
rect 440 480 455 500
rect 600 480 615 500
rect 760 480 775 500
rect 840 480 855 500
rect 925 480 940 500
rect 1120 480 1135 500
rect 40 180 55 438
rect 200 320 215 396
rect 175 310 215 320
rect 175 290 185 310
rect 205 290 215 310
rect 175 280 215 290
rect 15 170 55 180
rect 15 150 25 170
rect 45 150 55 170
rect 15 140 55 150
rect 40 4 55 140
rect 200 4 215 280
rect 280 273 295 396
rect 252 264 295 273
rect 252 237 261 264
rect 287 237 295 264
rect 252 230 295 237
rect 280 80 295 230
rect 440 131 455 438
rect 600 190 615 438
rect 570 180 615 190
rect 570 160 580 180
rect 600 160 615 180
rect 570 150 615 160
rect 410 121 455 131
rect 410 101 420 121
rect 440 101 455 121
rect 410 91 455 101
rect 280 70 320 80
rect 280 50 290 70
rect 310 50 320 70
rect 280 40 320 50
rect 280 4 295 40
rect 440 4 455 91
rect 600 4 615 150
rect 760 140 775 354
rect 840 223 855 354
rect 812 214 855 223
rect 812 187 821 214
rect 847 187 855 214
rect 812 180 855 187
rect 730 130 775 140
rect 730 110 740 130
rect 760 110 775 130
rect 730 100 775 110
rect 760 4 775 100
rect 840 4 855 180
rect 925 183 940 354
rect 1120 310 1135 438
rect 1095 300 1135 310
rect 1095 280 1105 300
rect 1125 280 1135 300
rect 1095 270 1135 280
rect 925 174 968 183
rect 925 147 934 174
rect 960 147 968 174
rect 925 140 968 147
rect 925 4 940 140
rect 1120 4 1135 270
rect 40 -100 55 -80
rect 200 -100 215 -80
rect 280 -100 295 -80
rect 440 -100 455 -80
rect 600 -100 615 -80
rect 760 -100 775 -80
rect 840 -100 855 -80
rect 925 -100 940 -80
rect 1120 -100 1135 -80
rect 340 -300 355 -280
rect 425 -300 440 -280
rect 600 -300 615 -280
rect 685 -300 700 -280
rect 860 -300 875 -280
rect 940 -300 955 -280
rect 1020 -300 1035 -280
rect 1100 -300 1115 -280
rect 340 -510 355 -384
rect 310 -524 355 -510
rect 310 -550 320 -524
rect 346 -550 355 -524
rect 310 -560 355 -550
rect 340 -832 355 -560
rect 425 -420 440 -384
rect 425 -430 465 -420
rect 425 -450 434 -430
rect 456 -450 465 -430
rect 425 -460 465 -450
rect 425 -832 440 -460
rect 600 -570 615 -384
rect 575 -580 615 -570
rect 575 -600 584 -580
rect 606 -600 615 -580
rect 575 -610 615 -600
rect 600 -832 615 -610
rect 685 -410 700 -384
rect 685 -420 725 -410
rect 685 -440 694 -420
rect 716 -440 725 -420
rect 685 -450 725 -440
rect 685 -832 700 -450
rect 860 -570 875 -384
rect 835 -580 875 -570
rect 835 -600 844 -580
rect 866 -600 875 -580
rect 835 -610 875 -600
rect 860 -748 875 -610
rect 940 -630 955 -384
rect 1020 -510 1035 -384
rect 990 -524 1035 -510
rect 990 -550 1000 -524
rect 1026 -550 1035 -524
rect 990 -560 1035 -550
rect 910 -644 955 -630
rect 910 -670 920 -644
rect 946 -670 955 -644
rect 910 -680 955 -670
rect 940 -748 955 -680
rect 1020 -748 1035 -560
rect 1100 -630 1115 -384
rect 1070 -644 1115 -630
rect 1070 -670 1080 -644
rect 1106 -670 1115 -644
rect 1070 -680 1115 -670
rect 1100 -748 1115 -680
rect 340 -936 355 -916
rect 425 -936 440 -916
rect 600 -936 615 -916
rect 685 -936 700 -916
rect 860 -936 875 -916
rect 940 -936 955 -916
rect 1020 -936 1035 -916
rect 1100 -936 1115 -916
rect 340 -1096 355 -1076
rect 425 -1096 440 -1076
rect 600 -1096 615 -1076
rect 685 -1096 700 -1076
rect 340 -1231 355 -1180
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1267 355 -1241
rect 310 -1281 355 -1267
rect 340 -1341 355 -1281
rect 310 -1351 355 -1341
rect 310 -1377 320 -1351
rect 346 -1377 355 -1351
rect 310 -1391 355 -1377
rect 340 -1517 355 -1391
rect 425 -1441 440 -1180
rect 600 -1371 615 -1180
rect 575 -1381 615 -1371
rect 575 -1401 584 -1381
rect 606 -1401 615 -1381
rect 575 -1411 615 -1401
rect 425 -1451 465 -1441
rect 425 -1471 434 -1451
rect 456 -1471 465 -1451
rect 425 -1481 465 -1471
rect 425 -1517 440 -1481
rect 600 -1517 615 -1411
rect 685 -1301 700 -1180
rect 685 -1311 725 -1301
rect 685 -1331 694 -1311
rect 716 -1331 725 -1311
rect 685 -1341 725 -1331
rect 685 -1517 700 -1341
rect 340 -1621 355 -1601
rect 425 -1621 440 -1601
rect 600 -1621 615 -1601
rect 685 -1621 700 -1601
rect 37 -1761 52 -1741
rect 197 -1761 212 -1741
rect 277 -1761 292 -1741
rect 437 -1761 452 -1741
rect 597 -1761 612 -1741
rect 790 -1761 805 -1741
rect 870 -1761 885 -1741
rect 955 -1761 970 -1741
rect 1150 -1761 1165 -1741
rect 37 -1981 52 -1845
rect 12 -1991 52 -1981
rect 12 -2011 22 -1991
rect 42 -2011 52 -1991
rect 12 -2021 52 -2011
rect 37 -2269 52 -2021
rect 197 -2121 212 -1845
rect 277 -1881 292 -1845
rect 277 -1891 317 -1881
rect 277 -1911 287 -1891
rect 307 -1911 317 -1891
rect 277 -1921 317 -1911
rect 277 -2071 292 -1921
rect 437 -1932 452 -1845
rect 407 -1942 452 -1932
rect 407 -1962 417 -1942
rect 437 -1962 452 -1942
rect 407 -1972 452 -1962
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2105 292 -2078
rect 249 -2114 292 -2105
rect 172 -2131 212 -2121
rect 172 -2151 182 -2131
rect 202 -2151 212 -2131
rect 172 -2161 212 -2151
rect 197 -2227 212 -2161
rect 277 -2227 292 -2114
rect 437 -2269 452 -1972
rect 597 -1991 612 -1845
rect 790 -1941 805 -1845
rect 760 -1951 805 -1941
rect 760 -1971 770 -1951
rect 790 -1971 805 -1951
rect 760 -1981 805 -1971
rect 567 -2001 612 -1991
rect 567 -2021 577 -2001
rect 597 -2021 612 -2001
rect 567 -2031 612 -2021
rect 597 -2269 612 -2031
rect 790 -2185 805 -1981
rect 870 -2021 885 -1845
rect 842 -2028 885 -2021
rect 842 -2055 851 -2028
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 870 -2185 885 -2064
rect 955 -1981 970 -1845
rect 955 -1988 998 -1981
rect 955 -2015 964 -1988
rect 990 -2015 998 -1988
rect 955 -2024 998 -2015
rect 955 -2185 970 -2024
rect 1150 -2111 1165 -1845
rect 1125 -2121 1165 -2111
rect 1125 -2141 1135 -2121
rect 1155 -2141 1165 -2121
rect 1125 -2151 1165 -2141
rect 1150 -2269 1165 -2151
rect 37 -2331 52 -2311
rect 197 -2331 212 -2311
rect 277 -2331 292 -2311
rect 437 -2331 452 -2311
rect 597 -2331 612 -2311
rect 790 -2331 805 -2311
rect 870 -2331 885 -2311
rect 955 -2331 970 -2311
rect 1150 -2331 1165 -2311
<< polycont >>
rect 185 290 205 310
rect 25 150 45 170
rect 261 237 287 264
rect 580 160 600 180
rect 420 101 440 121
rect 290 50 310 70
rect 821 187 847 214
rect 740 110 760 130
rect 1105 280 1125 300
rect 934 147 960 174
rect 320 -550 346 -524
rect 434 -450 456 -430
rect 584 -600 606 -580
rect 694 -440 716 -420
rect 844 -600 866 -580
rect 1000 -550 1026 -524
rect 920 -670 946 -644
rect 1080 -670 1106 -644
rect 320 -1267 346 -1241
rect 320 -1377 346 -1351
rect 584 -1401 606 -1381
rect 434 -1471 456 -1451
rect 694 -1331 716 -1311
rect 22 -2011 42 -1991
rect 287 -1911 307 -1891
rect 417 -1962 437 -1942
rect 258 -2105 284 -2078
rect 182 -2151 202 -2131
rect 770 -1971 790 -1951
rect 577 -2021 597 -2001
rect 851 -2055 877 -2028
rect 964 -2015 990 -1988
rect 1135 -2141 1155 -2121
<< locali >>
rect -70 590 1390 610
rect -70 550 -40 590
rect 0 550 40 590
rect 80 550 120 590
rect 160 550 200 590
rect 240 550 280 590
rect 320 550 360 590
rect 400 550 440 590
rect 480 550 520 590
rect 560 550 600 590
rect 640 550 680 590
rect 720 550 760 590
rect 800 550 840 590
rect 880 550 920 590
rect 960 550 1000 590
rect 1040 550 1080 590
rect 1120 550 1160 590
rect 1200 550 1240 590
rect 1280 550 1320 590
rect 1360 550 1390 590
rect -70 530 1390 550
rect -10 480 20 530
rect 150 480 180 530
rect 390 480 420 530
rect 550 480 580 530
rect 710 480 740 530
rect 1070 480 1100 530
rect 1310 490 1330 530
rect 1370 490 1390 530
rect -10 472 30 480
rect -10 448 -2 472
rect 22 448 30 472
rect -10 438 30 448
rect 70 472 110 480
rect 70 448 78 472
rect 102 448 110 472
rect 70 438 110 448
rect 80 310 110 438
rect 150 473 190 480
rect 150 405 158 473
rect 182 405 190 473
rect 150 396 190 405
rect 305 472 345 480
rect 305 404 313 472
rect 337 404 345 472
rect 390 472 430 480
rect 390 448 398 472
rect 422 448 430 472
rect 390 438 430 448
rect 470 472 510 480
rect 470 448 478 472
rect 502 448 510 472
rect 470 438 510 448
rect 550 472 590 480
rect 550 448 558 472
rect 582 448 590 472
rect 550 438 590 448
rect 630 472 670 480
rect 630 448 638 472
rect 662 448 670 472
rect 630 438 670 448
rect 305 396 345 404
rect 175 310 215 320
rect 80 290 185 310
rect 205 290 215 310
rect 80 280 215 290
rect 15 170 55 180
rect -30 150 25 170
rect 45 150 55 170
rect -30 140 55 150
rect 80 4 110 280
rect 252 264 295 273
rect 252 237 261 264
rect 287 237 295 264
rect 252 230 295 237
rect 315 131 345 396
rect 480 180 510 438
rect 570 180 610 190
rect 480 160 580 180
rect 600 160 610 180
rect 480 150 610 160
rect 231 121 450 131
rect 231 101 420 121
rect 440 101 450 121
rect 231 4 261 101
rect 410 91 450 101
rect 280 70 320 80
rect 280 50 290 70
rect 310 50 320 70
rect 280 40 320 50
rect 480 4 510 150
rect 640 130 670 438
rect 710 452 750 480
rect 710 384 718 452
rect 742 384 750 452
rect 710 354 750 384
rect 950 445 990 480
rect 950 377 958 445
rect 982 377 990 445
rect 1070 472 1110 480
rect 1070 448 1078 472
rect 1102 448 1110 472
rect 1070 438 1110 448
rect 1150 472 1190 480
rect 1150 448 1158 472
rect 1182 448 1190 472
rect 1150 438 1190 448
rect 950 354 990 377
rect 950 310 980 354
rect 874 300 1135 310
rect 874 280 1105 300
rect 1125 280 1135 300
rect 700 273 740 280
rect 700 247 707 273
rect 733 270 740 273
rect 874 270 904 280
rect 1095 270 1135 280
rect 733 247 904 270
rect 700 240 904 247
rect 812 214 855 223
rect 812 187 821 214
rect 847 187 855 214
rect 812 180 855 187
rect 730 130 770 140
rect 640 110 740 130
rect 760 110 770 130
rect 640 100 770 110
rect 640 4 670 100
rect 790 70 830 80
rect 874 70 904 240
rect 925 174 968 183
rect 925 147 934 174
rect 960 147 968 174
rect 925 140 968 147
rect 1160 120 1190 438
rect 1310 450 1390 490
rect 1310 310 1330 450
rect 1370 310 1390 450
rect 1310 270 1390 310
rect 1310 230 1330 270
rect 1370 230 1390 270
rect 1310 190 1390 230
rect 1310 150 1330 190
rect 1370 150 1390 190
rect 1160 90 1230 120
rect 1310 110 1390 150
rect 790 50 800 70
rect 820 50 990 70
rect 790 40 990 50
rect 793 4 823 40
rect 960 4 990 40
rect 1160 4 1190 90
rect -10 -20 30 4
rect -10 -60 -4 -20
rect 26 -60 30 -20
rect -10 -80 30 -60
rect 70 -20 110 4
rect 70 -60 73 -20
rect 103 -60 110 -20
rect 70 -80 110 -60
rect 150 -20 190 4
rect 150 -60 156 -20
rect 186 -60 190 -20
rect 150 -80 190 -60
rect 227 -20 267 4
rect 227 -60 232 -20
rect 262 -60 267 -20
rect 227 -80 267 -60
rect 305 -20 345 4
rect 305 -60 310 -20
rect 340 -60 345 -20
rect 305 -80 345 -60
rect -10 -120 20 -80
rect 150 -120 180 -80
rect 315 -120 345 -80
rect 390 -20 430 4
rect 390 -60 396 -20
rect 426 -60 430 -20
rect 390 -80 430 -60
rect 470 -20 510 4
rect 470 -60 473 -20
rect 503 -60 510 -20
rect 470 -80 510 -60
rect 550 -20 590 4
rect 550 -60 556 -20
rect 586 -60 590 -20
rect 550 -80 590 -60
rect 630 -20 670 4
rect 630 -60 633 -20
rect 663 -60 670 -20
rect 630 -80 670 -60
rect 710 -20 750 4
rect 710 -60 716 -20
rect 746 -60 750 -20
rect 710 -80 750 -60
rect 788 -20 828 4
rect 788 -60 794 -20
rect 824 -60 828 -20
rect 788 -80 828 -60
rect 870 -20 910 4
rect 870 -60 876 -20
rect 906 -60 910 -20
rect 870 -80 910 -60
rect 950 -20 990 4
rect 950 -60 955 -20
rect 985 -60 990 -20
rect 950 -80 990 -60
rect 1070 -20 1110 4
rect 1070 -60 1076 -20
rect 1106 -60 1110 -20
rect 1070 -80 1110 -60
rect 1150 -20 1190 4
rect 1150 -60 1153 -20
rect 1183 -60 1190 -20
rect 1150 -80 1190 -60
rect 1310 70 1330 110
rect 1370 70 1390 110
rect 1310 30 1390 70
rect 1310 -10 1330 30
rect 1370 -10 1390 30
rect 1310 -50 1390 -10
rect 390 -120 420 -80
rect 550 -120 580 -80
rect 710 -120 740 -80
rect 870 -120 900 -80
rect 1070 -120 1100 -80
rect 1310 -90 1330 -50
rect 1370 -90 1390 -50
rect -130 -140 1245 -120
rect -130 -180 -50 -140
rect -10 -180 20 -140
rect 60 -180 90 -140
rect 130 -180 160 -140
rect 200 -180 310 -140
rect 350 -180 740 -140
rect 780 -180 800 -140
rect 840 -180 870 -140
rect 910 -180 940 -140
rect 980 -180 1100 -140
rect 1140 -180 1160 -140
rect 1200 -180 1245 -140
rect -130 -200 1245 -180
rect 1310 -130 1390 -90
rect 1310 -170 1330 -130
rect 1370 -170 1390 -130
rect -130 -1641 -50 -200
rect 290 -300 320 -200
rect 460 -300 490 -200
rect 290 -320 330 -300
rect 290 -360 296 -320
rect 326 -360 330 -320
rect 290 -384 330 -360
rect 370 -320 410 -300
rect 370 -360 375 -320
rect 405 -360 410 -320
rect 370 -384 410 -360
rect 450 -320 490 -300
rect 450 -360 453 -320
rect 483 -360 490 -320
rect 450 -384 490 -360
rect 550 -300 580 -200
rect 720 -300 750 -200
rect 550 -320 590 -300
rect 550 -360 556 -320
rect 586 -360 590 -320
rect 550 -384 590 -360
rect 630 -320 670 -300
rect 630 -360 635 -320
rect 665 -360 670 -320
rect 630 -384 670 -360
rect 710 -320 750 -300
rect 710 -360 713 -320
rect 743 -360 750 -320
rect 710 -384 750 -360
rect 810 -300 840 -200
rect 970 -300 1000 -200
rect 1130 -300 1160 -200
rect 1310 -210 1390 -170
rect 1310 -250 1330 -210
rect 1370 -250 1390 -210
rect 1310 -290 1390 -250
rect 810 -319 850 -300
rect 810 -359 816 -319
rect 846 -359 850 -319
rect 810 -384 850 -359
rect 890 -320 930 -300
rect 890 -360 895 -320
rect 925 -360 930 -320
rect 890 -384 930 -360
rect 970 -319 1010 -300
rect 970 -359 976 -319
rect 1006 -359 1010 -319
rect 970 -384 1010 -359
rect 1050 -319 1090 -300
rect 1050 -359 1056 -319
rect 1086 -359 1090 -319
rect 1050 -384 1090 -359
rect 1130 -319 1170 -300
rect 1130 -359 1136 -319
rect 1166 -359 1170 -319
rect 1130 -384 1170 -359
rect 1310 -330 1330 -290
rect 1370 -330 1390 -290
rect 1310 -370 1390 -330
rect 374 -480 404 -384
rect 634 -420 664 -384
rect 425 -430 664 -420
rect 425 -450 434 -430
rect 456 -450 664 -430
rect 685 -420 725 -410
rect 890 -420 920 -384
rect 1060 -420 1090 -384
rect 685 -440 694 -420
rect 716 -440 1090 -420
rect 685 -450 1090 -440
rect 425 -460 465 -450
rect 634 -470 664 -450
rect 374 -510 490 -480
rect 634 -500 750 -470
rect 310 -524 355 -510
rect 310 -550 320 -524
rect 346 -550 355 -524
rect 310 -560 355 -550
rect 460 -580 490 -510
rect 575 -580 615 -570
rect 460 -600 584 -580
rect 606 -600 615 -580
rect 460 -610 615 -600
rect 460 -832 490 -610
rect 720 -832 750 -500
rect 990 -524 1035 -510
rect 990 -550 1000 -524
rect 1026 -550 1035 -524
rect 990 -560 1035 -550
rect 1060 -560 1090 -450
rect 1310 -410 1330 -370
rect 1370 -410 1390 -370
rect 1310 -450 1390 -410
rect 1310 -490 1330 -450
rect 1370 -490 1390 -450
rect 1310 -530 1390 -490
rect 835 -580 875 -570
rect 835 -600 844 -580
rect 866 -600 875 -580
rect 1060 -590 1170 -560
rect 835 -610 875 -600
rect 910 -644 955 -630
rect 910 -670 920 -644
rect 946 -670 955 -644
rect 910 -680 955 -670
rect 1070 -644 1115 -630
rect 1070 -670 1080 -644
rect 1106 -670 1115 -644
rect 1070 -680 1115 -670
rect 1140 -748 1170 -590
rect 1310 -570 1330 -530
rect 1370 -570 1390 -530
rect 1310 -610 1390 -570
rect 1310 -650 1330 -610
rect 1370 -650 1390 -610
rect 1310 -690 1390 -650
rect 290 -840 330 -832
rect 290 -908 298 -840
rect 322 -908 330 -840
rect 290 -916 330 -908
rect 450 -840 490 -832
rect 450 -908 458 -840
rect 482 -908 490 -840
rect 450 -916 490 -908
rect 550 -840 590 -832
rect 550 -908 558 -840
rect 582 -908 590 -840
rect 550 -916 590 -908
rect 710 -840 750 -832
rect 710 -908 718 -840
rect 742 -908 750 -840
rect 710 -916 750 -908
rect 810 -780 850 -748
rect 810 -899 818 -780
rect 841 -899 850 -780
rect 810 -916 850 -899
rect 1129 -776 1171 -748
rect 1129 -897 1137 -776
rect 1163 -897 1171 -776
rect 290 -966 320 -916
rect 550 -966 580 -916
rect 810 -966 840 -916
rect 1129 -917 1171 -897
rect 1310 -886 1330 -690
rect 1370 -886 1390 -690
rect 1310 -926 1390 -886
rect 1310 -966 1330 -926
rect 1370 -966 1390 -926
rect 280 -986 1390 -966
rect 280 -1026 310 -986
rect 350 -1026 390 -986
rect 430 -1026 830 -986
rect 870 -1026 910 -986
rect 950 -1026 990 -986
rect 1030 -1026 1070 -986
rect 1110 -1026 1270 -986
rect 1310 -1006 1390 -986
rect 1310 -1026 1330 -1006
rect 280 -1046 1330 -1026
rect 1370 -1046 1390 -1006
rect 290 -1096 320 -1046
rect 290 -1104 330 -1096
rect 290 -1172 298 -1104
rect 322 -1172 330 -1104
rect 290 -1180 330 -1172
rect 450 -1104 492 -1094
rect 450 -1172 458 -1104
rect 484 -1172 492 -1104
rect 450 -1180 492 -1172
rect 550 -1096 580 -1046
rect 1310 -1086 1390 -1046
rect 550 -1104 590 -1096
rect 550 -1172 558 -1104
rect 582 -1172 590 -1104
rect 550 -1180 590 -1172
rect 710 -1104 750 -1096
rect 710 -1172 718 -1104
rect 742 -1172 750 -1104
rect 1128 -1112 1170 -1105
rect 1128 -1138 1136 -1112
rect 1162 -1138 1170 -1112
rect 1128 -1146 1170 -1138
rect 710 -1180 750 -1172
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1267 355 -1241
rect 310 -1281 355 -1267
rect 310 -1351 355 -1341
rect 310 -1377 320 -1351
rect 346 -1377 355 -1351
rect 460 -1371 490 -1180
rect 720 -1201 750 -1180
rect 634 -1231 750 -1201
rect 310 -1391 355 -1377
rect 374 -1381 615 -1371
rect 374 -1401 584 -1381
rect 606 -1401 615 -1381
rect 374 -1517 404 -1401
rect 575 -1411 615 -1401
rect 425 -1451 465 -1441
rect 634 -1451 664 -1231
rect 1140 -1301 1170 -1146
rect 685 -1311 1170 -1301
rect 685 -1331 694 -1311
rect 716 -1331 1170 -1311
rect 1310 -1126 1330 -1086
rect 1370 -1126 1390 -1086
rect 1310 -1211 1390 -1126
rect 1310 -1251 1330 -1211
rect 1370 -1251 1390 -1211
rect 1310 -1291 1390 -1251
rect 1310 -1331 1330 -1291
rect 1370 -1331 1390 -1291
rect 685 -1341 725 -1331
rect 1053 -1420 1083 -1331
rect 1310 -1371 1390 -1331
rect 1310 -1411 1330 -1371
rect 1370 -1411 1390 -1371
rect 425 -1471 434 -1451
rect 456 -1471 664 -1451
rect 1043 -1427 1085 -1420
rect 1043 -1453 1051 -1427
rect 1077 -1453 1085 -1427
rect 1043 -1461 1085 -1453
rect 1310 -1451 1390 -1411
rect 425 -1481 664 -1471
rect 634 -1517 664 -1481
rect 1310 -1491 1330 -1451
rect 1370 -1491 1390 -1451
rect 290 -1541 330 -1517
rect 290 -1581 296 -1541
rect 326 -1581 330 -1541
rect 290 -1601 330 -1581
rect 370 -1541 410 -1517
rect 370 -1581 375 -1541
rect 405 -1581 410 -1541
rect 370 -1601 410 -1581
rect 450 -1541 490 -1517
rect 450 -1581 453 -1541
rect 483 -1581 490 -1541
rect 450 -1601 490 -1581
rect 290 -1641 320 -1601
rect 460 -1641 490 -1601
rect 550 -1541 590 -1517
rect 550 -1581 556 -1541
rect 586 -1581 590 -1541
rect 550 -1601 590 -1581
rect 630 -1541 670 -1517
rect 630 -1581 635 -1541
rect 665 -1581 670 -1541
rect 630 -1601 670 -1581
rect 710 -1541 750 -1517
rect 710 -1581 713 -1541
rect 743 -1581 750 -1541
rect 710 -1601 750 -1581
rect 550 -1641 580 -1601
rect 720 -1641 750 -1601
rect 1310 -1531 1390 -1491
rect 1310 -1571 1330 -1531
rect 1370 -1571 1390 -1531
rect 1310 -1611 1390 -1571
rect -130 -1661 1250 -1641
rect -130 -1701 -70 -1661
rect -30 -1701 0 -1661
rect 40 -1701 70 -1661
rect 110 -1701 140 -1661
rect 180 -1701 300 -1661
rect 340 -1701 750 -1661
rect 790 -1701 820 -1661
rect 860 -1701 890 -1661
rect 930 -1701 960 -1661
rect 1000 -1701 1100 -1661
rect 1140 -1701 1170 -1661
rect 1210 -1701 1250 -1661
rect -130 -1721 1250 -1701
rect 1310 -1651 1330 -1611
rect 1370 -1651 1390 -1611
rect 1310 -1691 1390 -1651
rect -13 -1761 17 -1721
rect 147 -1761 177 -1721
rect 312 -1761 342 -1721
rect -13 -1781 27 -1761
rect -13 -1821 -7 -1781
rect 23 -1821 27 -1781
rect -13 -1845 27 -1821
rect 67 -1781 107 -1761
rect 67 -1821 70 -1781
rect 100 -1821 107 -1781
rect 67 -1845 107 -1821
rect 147 -1781 187 -1761
rect 147 -1821 153 -1781
rect 183 -1821 187 -1781
rect 147 -1845 187 -1821
rect 224 -1781 264 -1761
rect 224 -1821 229 -1781
rect 259 -1821 264 -1781
rect 224 -1845 264 -1821
rect 302 -1781 342 -1761
rect 302 -1821 307 -1781
rect 337 -1821 342 -1781
rect 302 -1845 342 -1821
rect 387 -1761 417 -1721
rect 547 -1761 577 -1721
rect 740 -1761 770 -1721
rect 900 -1761 930 -1721
rect 1100 -1761 1130 -1721
rect 1310 -1731 1330 -1691
rect 1370 -1731 1390 -1691
rect 387 -1781 427 -1761
rect 387 -1821 393 -1781
rect 423 -1821 427 -1781
rect 387 -1845 427 -1821
rect 467 -1781 507 -1761
rect 467 -1821 470 -1781
rect 500 -1821 507 -1781
rect 467 -1845 507 -1821
rect 547 -1781 587 -1761
rect 547 -1821 553 -1781
rect 583 -1821 587 -1781
rect 547 -1845 587 -1821
rect 627 -1781 667 -1761
rect 627 -1821 630 -1781
rect 660 -1821 667 -1781
rect 627 -1845 667 -1821
rect 740 -1781 780 -1761
rect 740 -1821 745 -1781
rect 776 -1821 780 -1781
rect 740 -1845 780 -1821
rect 818 -1781 858 -1761
rect 818 -1821 824 -1781
rect 854 -1821 858 -1781
rect 818 -1845 858 -1821
rect 900 -1781 940 -1761
rect 900 -1821 906 -1781
rect 936 -1821 940 -1781
rect 900 -1845 940 -1821
rect 980 -1781 1020 -1761
rect 980 -1821 985 -1781
rect 1015 -1821 1020 -1781
rect 980 -1845 1020 -1821
rect 1100 -1781 1140 -1761
rect 1100 -1821 1106 -1781
rect 1136 -1821 1140 -1781
rect 1100 -1845 1140 -1821
rect 1180 -1781 1220 -1761
rect 1180 -1821 1183 -1781
rect 1213 -1821 1220 -1781
rect 1180 -1845 1220 -1821
rect 12 -1991 52 -1981
rect -30 -2011 22 -1991
rect 42 -2011 52 -1991
rect -30 -2021 52 -2011
rect 77 -2121 107 -1845
rect 228 -1942 258 -1845
rect 277 -1891 317 -1881
rect 277 -1911 287 -1891
rect 307 -1911 317 -1891
rect 277 -1921 317 -1911
rect 407 -1942 447 -1932
rect 228 -1962 417 -1942
rect 437 -1962 447 -1942
rect 228 -1972 447 -1962
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2105 292 -2078
rect 249 -2114 292 -2105
rect 77 -2131 212 -2121
rect 77 -2151 182 -2131
rect 202 -2151 212 -2131
rect 77 -2269 107 -2151
rect 172 -2161 212 -2151
rect 312 -2227 342 -1972
rect -13 -2279 27 -2269
rect -13 -2303 -5 -2279
rect 19 -2303 27 -2279
rect -13 -2311 27 -2303
rect 67 -2279 107 -2269
rect 67 -2303 75 -2279
rect 99 -2303 107 -2279
rect 67 -2311 107 -2303
rect 147 -2235 187 -2227
rect 147 -2303 155 -2235
rect 179 -2303 187 -2235
rect 147 -2311 187 -2303
rect 302 -2235 342 -2227
rect 302 -2303 311 -2235
rect 335 -2303 342 -2235
rect 477 -1991 507 -1845
rect 637 -1941 667 -1845
rect 823 -1881 853 -1845
rect 990 -1881 1020 -1845
rect 820 -1891 1020 -1881
rect 820 -1911 830 -1891
rect 850 -1911 1020 -1891
rect 820 -1921 860 -1911
rect 637 -1951 800 -1941
rect 637 -1971 770 -1951
rect 790 -1971 800 -1951
rect 477 -2001 607 -1991
rect 477 -2021 577 -2001
rect 597 -2021 607 -2001
rect 477 -2269 507 -2021
rect 567 -2031 607 -2021
rect 637 -2269 667 -1971
rect 760 -1981 800 -1971
rect 842 -2028 885 -2021
rect 842 -2055 851 -2028
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 904 -2081 934 -1911
rect 1190 -1931 1220 -1845
rect 1310 -1771 1390 -1731
rect 1310 -1811 1330 -1771
rect 1370 -1811 1390 -1771
rect 1310 -1851 1390 -1811
rect 1310 -1891 1330 -1851
rect 1370 -1891 1390 -1851
rect 1310 -1931 1390 -1891
rect 1190 -1961 1260 -1931
rect 955 -1988 998 -1981
rect 955 -2015 964 -1988
rect 990 -2015 998 -1988
rect 955 -2024 998 -2015
rect 730 -2088 934 -2081
rect 730 -2114 737 -2088
rect 763 -2111 934 -2088
rect 763 -2114 770 -2111
rect 730 -2121 770 -2114
rect 904 -2121 934 -2111
rect 1125 -2121 1165 -2111
rect 904 -2141 1135 -2121
rect 1155 -2141 1165 -2121
rect 904 -2151 1165 -2141
rect 980 -2185 1010 -2151
rect 302 -2311 342 -2303
rect 387 -2279 427 -2269
rect 387 -2303 395 -2279
rect 419 -2303 427 -2279
rect 387 -2311 427 -2303
rect 467 -2279 507 -2269
rect 467 -2303 475 -2279
rect 499 -2303 507 -2279
rect 467 -2311 507 -2303
rect 547 -2279 587 -2269
rect 547 -2303 555 -2279
rect 579 -2303 587 -2279
rect 547 -2311 587 -2303
rect 627 -2279 667 -2269
rect 627 -2303 635 -2279
rect 659 -2303 667 -2279
rect 627 -2311 667 -2303
rect 740 -2221 780 -2185
rect 740 -2289 748 -2221
rect 772 -2289 780 -2221
rect 740 -2311 780 -2289
rect 980 -2212 1020 -2185
rect 980 -2280 988 -2212
rect 1012 -2280 1020 -2212
rect 1190 -2269 1220 -1961
rect 980 -2311 1020 -2280
rect 1100 -2279 1140 -2269
rect 1100 -2303 1108 -2279
rect 1132 -2303 1140 -2279
rect 1100 -2311 1140 -2303
rect 1180 -2279 1220 -2269
rect 1180 -2303 1188 -2279
rect 1212 -2303 1220 -2279
rect 1180 -2311 1220 -2303
rect 1310 -1971 1330 -1931
rect 1370 -1971 1390 -1931
rect 1310 -2011 1390 -1971
rect 1310 -2051 1330 -2011
rect 1370 -2051 1390 -2011
rect 1310 -2091 1390 -2051
rect 1310 -2131 1330 -2091
rect 1370 -2131 1390 -2091
rect 1310 -2261 1390 -2131
rect 1310 -2301 1330 -2261
rect 1370 -2301 1390 -2261
rect -13 -2361 17 -2311
rect 147 -2361 177 -2311
rect 387 -2361 417 -2311
rect 547 -2361 577 -2311
rect 740 -2361 770 -2311
rect 1100 -2361 1130 -2311
rect 1310 -2361 1390 -2301
rect -73 -2371 1390 -2361
rect -73 -2381 1330 -2371
rect -73 -2421 -40 -2381
rect 0 -2421 40 -2381
rect 80 -2421 120 -2381
rect 160 -2421 200 -2381
rect 240 -2421 280 -2381
rect 320 -2421 360 -2381
rect 400 -2421 440 -2381
rect 480 -2421 520 -2381
rect 560 -2421 600 -2381
rect 640 -2421 680 -2381
rect 720 -2421 760 -2381
rect 800 -2421 840 -2381
rect 880 -2421 920 -2381
rect 960 -2421 1000 -2381
rect 1040 -2421 1080 -2381
rect 1120 -2421 1160 -2381
rect 1200 -2421 1240 -2381
rect 1280 -2411 1330 -2381
rect 1370 -2411 1390 -2371
rect 1280 -2421 1390 -2411
rect -73 -2441 1390 -2421
<< viali >>
rect 261 237 287 264
rect 290 50 310 70
rect 707 247 733 273
rect 821 187 847 214
rect 934 147 960 174
rect 800 50 820 70
rect 232 -60 262 -20
rect 375 -360 405 -320
rect 1056 -359 1086 -319
rect 320 -550 346 -524
rect 584 -600 606 -580
rect 1000 -550 1026 -524
rect 844 -600 866 -580
rect 920 -670 946 -644
rect 1080 -670 1106 -644
rect 1137 -897 1163 -776
rect 458 -1172 484 -1104
rect 1136 -1138 1162 -1112
rect 320 -1267 346 -1241
rect 320 -1377 346 -1351
rect 584 -1401 606 -1381
rect 1051 -1453 1077 -1427
rect 375 -1581 405 -1541
rect 229 -1821 259 -1781
rect 287 -1911 307 -1891
rect 258 -2105 284 -2078
rect 830 -1911 850 -1891
rect 851 -2055 877 -2028
rect 964 -2015 990 -1988
rect 737 -2114 763 -2088
<< metal1 >>
rect 700 273 740 280
rect 252 264 295 273
rect 252 237 261 264
rect 287 237 295 264
rect 700 247 707 273
rect 733 247 740 273
rect 700 240 740 247
rect 252 230 295 237
rect 812 214 855 223
rect 812 187 821 214
rect 847 187 855 214
rect 812 180 855 187
rect 925 174 968 183
rect 925 147 934 174
rect 960 147 968 174
rect 925 140 968 147
rect 280 70 320 80
rect 790 70 830 80
rect 280 50 290 70
rect 310 50 800 70
rect 820 50 830 70
rect 280 40 830 50
rect 227 -20 267 4
rect 227 -60 232 -20
rect 262 -60 267 -20
rect 227 -80 267 -60
rect 370 -320 410 -300
rect 370 -360 375 -320
rect 405 -360 410 -320
rect 370 -384 410 -360
rect 1050 -319 1090 -300
rect 1050 -359 1056 -319
rect 1086 -359 1090 -319
rect 1050 -384 1090 -359
rect 310 -524 355 -510
rect 310 -550 320 -524
rect 346 -550 355 -524
rect 310 -560 355 -550
rect 990 -524 1035 -510
rect 990 -550 1000 -524
rect 1026 -550 1035 -524
rect 990 -560 1035 -550
rect 575 -580 615 -570
rect 835 -580 875 -570
rect 575 -600 584 -580
rect 606 -600 844 -580
rect 866 -600 875 -580
rect 575 -610 875 -600
rect 910 -644 955 -630
rect 910 -670 920 -644
rect 946 -670 955 -644
rect 910 -680 955 -670
rect 1070 -644 1115 -630
rect 1070 -670 1080 -644
rect 1106 -670 1115 -644
rect 1070 -680 1115 -670
rect 1129 -776 1171 -748
rect 1129 -897 1137 -776
rect 1163 -897 1171 -776
rect 1129 -917 1171 -897
rect 450 -1104 492 -1094
rect 450 -1172 458 -1104
rect 484 -1172 492 -1104
rect 1128 -1112 1170 -1105
rect 1128 -1138 1136 -1112
rect 1162 -1138 1170 -1112
rect 1128 -1146 1170 -1138
rect 450 -1180 492 -1172
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1267 355 -1241
rect 310 -1281 355 -1267
rect 310 -1351 355 -1341
rect 310 -1377 320 -1351
rect 346 -1377 355 -1351
rect 310 -1391 355 -1377
rect 575 -1381 615 -1371
rect 575 -1401 584 -1381
rect 606 -1401 615 -1381
rect 575 -1411 615 -1401
rect 1043 -1427 1085 -1420
rect 1043 -1453 1051 -1427
rect 1077 -1453 1085 -1427
rect 1043 -1461 1085 -1453
rect 370 -1541 410 -1517
rect 370 -1581 375 -1541
rect 405 -1581 410 -1541
rect 370 -1601 410 -1581
rect 224 -1781 264 -1761
rect 224 -1821 229 -1781
rect 259 -1821 264 -1781
rect 224 -1845 264 -1821
rect 277 -1891 860 -1881
rect 277 -1911 287 -1891
rect 307 -1911 830 -1891
rect 850 -1911 860 -1891
rect 277 -1921 317 -1911
rect 820 -1921 860 -1911
rect 955 -1988 998 -1981
rect 955 -2015 964 -1988
rect 990 -2015 998 -1988
rect 842 -2028 885 -2021
rect 955 -2024 998 -2015
rect 842 -2055 851 -2028
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2105 292 -2078
rect 249 -2114 292 -2105
rect 730 -2088 770 -2081
rect 730 -2114 737 -2088
rect 763 -2114 770 -2088
rect 730 -2121 770 -2114
<< via1 >>
rect 261 237 287 264
rect 707 247 733 273
rect 821 187 847 214
rect 934 147 960 174
rect 232 -60 262 -20
rect 375 -360 405 -320
rect 1056 -359 1086 -319
rect 320 -550 346 -524
rect 1000 -550 1026 -524
rect 920 -670 946 -644
rect 1080 -670 1106 -644
rect 1137 -897 1163 -776
rect 458 -1172 484 -1104
rect 1136 -1138 1162 -1112
rect 320 -1267 346 -1241
rect 320 -1377 346 -1351
rect 1051 -1453 1077 -1427
rect 375 -1581 405 -1541
rect 229 -1821 259 -1781
rect 964 -2015 990 -1988
rect 851 -2055 877 -2028
rect 258 -2105 284 -2078
rect 737 -2114 763 -2088
<< metal2 >>
rect 700 273 740 280
rect 252 264 707 273
rect 252 237 261 264
rect 287 247 707 264
rect 733 247 740 273
rect 287 243 740 247
rect 287 237 295 243
rect 700 240 740 243
rect 252 230 295 237
rect 812 214 855 223
rect 812 210 821 214
rect 690 187 821 210
rect 847 187 855 214
rect 690 180 855 187
rect 227 -20 267 4
rect 227 -60 232 -20
rect 262 -60 267 -20
rect 227 -80 267 -60
rect 230 -520 260 -80
rect 690 -140 720 180
rect 925 174 968 183
rect 925 147 934 174
rect 960 170 968 174
rect 960 147 1040 170
rect 925 140 1040 147
rect 375 -170 720 -140
rect 1010 -140 1040 140
rect 1010 -170 1080 -140
rect 375 -300 405 -170
rect 1050 -300 1080 -170
rect 370 -320 410 -300
rect 370 -360 375 -320
rect 405 -360 410 -320
rect 370 -384 410 -360
rect 1050 -319 1090 -300
rect 1050 -359 1056 -319
rect 1086 -359 1090 -319
rect 1050 -384 1090 -359
rect 310 -520 355 -510
rect 990 -520 1035 -510
rect 230 -524 1035 -520
rect 230 -550 320 -524
rect 346 -550 1000 -524
rect 1026 -550 1035 -524
rect 310 -560 355 -550
rect 990 -560 1035 -550
rect 910 -644 955 -630
rect 910 -650 920 -644
rect 770 -670 920 -650
rect 946 -670 955 -644
rect 770 -680 955 -670
rect 1070 -644 1240 -630
rect 1070 -670 1080 -644
rect 1106 -660 1240 -644
rect 1106 -670 1115 -660
rect 1070 -680 1115 -670
rect 770 -986 800 -680
rect 462 -1016 800 -986
rect 1129 -776 1171 -748
rect 1129 -897 1137 -776
rect 1163 -897 1171 -776
rect 1129 -917 1171 -897
rect 462 -1094 492 -1016
rect 450 -1104 492 -1094
rect 450 -1172 458 -1104
rect 484 -1172 492 -1104
rect 1129 -1105 1159 -917
rect 1128 -1112 1170 -1105
rect 1128 -1138 1136 -1112
rect 1162 -1138 1170 -1112
rect 1128 -1146 1170 -1138
rect 450 -1180 492 -1172
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1251 355 -1241
rect 1210 -1251 1240 -660
rect 346 -1267 1240 -1251
rect 310 -1281 1240 -1267
rect 310 -1351 355 -1341
rect 227 -1377 320 -1351
rect 346 -1377 355 -1351
rect 227 -1381 355 -1377
rect 227 -1761 257 -1381
rect 310 -1391 355 -1381
rect 1043 -1427 1085 -1420
rect 1043 -1453 1051 -1427
rect 1077 -1453 1085 -1427
rect 1043 -1461 1085 -1453
rect 370 -1541 410 -1517
rect 370 -1581 375 -1541
rect 405 -1581 410 -1541
rect 370 -1601 410 -1581
rect 375 -1671 405 -1601
rect 375 -1701 720 -1671
rect 224 -1781 264 -1761
rect 224 -1821 229 -1781
rect 259 -1821 264 -1781
rect 224 -1845 264 -1821
rect 690 -2021 720 -1701
rect 1050 -1981 1080 -1461
rect 955 -1988 1080 -1981
rect 955 -2015 964 -1988
rect 990 -2011 1080 -1988
rect 990 -2015 998 -2011
rect 690 -2028 885 -2021
rect 955 -2024 998 -2015
rect 690 -2051 851 -2028
rect 842 -2055 851 -2051
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2084 292 -2078
rect 730 -2084 770 -2081
rect 284 -2088 770 -2084
rect 284 -2105 737 -2088
rect 249 -2114 737 -2105
rect 763 -2114 770 -2088
rect 730 -2121 770 -2114
<< labels >>
rlabel locali 1200 100 1220 110 1 up
rlabel locali -20 150 0 160 1 fin
rlabel locali 1230 -1951 1250 -1941 1 dn
rlabel locali -20 -2011 0 -2001 1 fvco_8
rlabel locali 1340 -996 1360 -986 1 gnd!
rlabel locali -100 -906 -80 -886 1 vdd
<< end >>
