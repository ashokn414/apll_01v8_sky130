* NGSPICE file created from freq_div_2.ext - technology: sky130A


* Top level circuit freq_div_2

X0 q a_404_n776# vdd vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X1 a_239_n520# a_90_n776# a_835_n776# vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X2 a_404_n776# clk a_284_n776# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_517_n776# clk a_404_n776# vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X4 a_835_n776# a_284_n776# gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_517_n776# q gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_239_n520# clk a_517_n776# vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X7 q a_404_n776# gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_517_n776# a_90_n776# a_404_n776# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_239_n520# clk a_835_n776# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_90_n776# clk vdd vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X11 a_284_n776# a_239_n520# vdd vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X12 a_239_n520# a_90_n776# a_517_n776# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_404_n776# a_90_n776# a_284_n776# vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X14 a_90_n776# clk gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_835_n776# a_284_n776# vdd vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
X16 a_284_n776# a_239_n520# gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_517_n776# q vdd vdd sky130_fd_pr__pfet_01v8 w=1.3e+06u l=150000u
.end

