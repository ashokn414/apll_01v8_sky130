***cs_inverter circuit***
.param L=0.15
.param W=0.42
.include "/home/ashok/sky130_fd_pr/models/corners/tt.spice"
.include "sky130_fd_pr/models/r+c/res_typical__cap_typical__lin.spice"
.include "sky130_fd_pr/models/r+c/res_typical__cap_typical.spice"



***Netlist Description***
X1 N003 Vn 0 0 sky130_fd_pr__nfet_01v8 l={L} w={2*W}
X4 N002 Vp N001 VDD sky130_fd_pr__pfet_01v8 l={L} w={4*W}
X3 Out In N002 VDD sky130_fd_pr__pfet_01v8 l={L} w={4*W}
X2 Out In N003 0 sky130_fd_pr__nfet_01v8 l={L} w={2*W}
C1 Out 0 1f
V1 N001 0 1.8

***simulation commands***
vdd VDD 0 1.8
vp1 Vp 0 1.8 
vn1 Vn 0 -1.8
Vin2 In 0 0 pulse(0 1.8 0 10p 10p 0.5n 1n) 

.op
.tran 10p 6n
.end
