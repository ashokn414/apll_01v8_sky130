magic
tech sky130A
timestamp 1605504292
<< nwell >>
rect -65 -262 1480 300
<< nmos >>
rect 75 -776 90 -734
rect 269 -776 284 -734
rect 389 -776 404 -734
rect 502 -776 517 -734
rect 612 -776 627 -734
rect 820 -776 835 -734
rect 940 -776 955 -734
rect 1131 -776 1146 -734
rect 1320 -776 1335 -734
<< pmos >>
rect 75 -200 90 -70
rect 269 -200 284 -70
rect 389 -200 404 -70
rect 502 -200 517 -70
rect 612 -200 627 -70
rect 820 -200 835 -70
rect 940 -200 955 -70
rect 1131 -200 1146 -70
rect 1320 -200 1335 -70
<< ndiff >>
rect 5 -744 75 -734
rect 5 -764 15 -744
rect 45 -764 75 -744
rect 5 -776 75 -764
rect 90 -744 159 -734
rect 90 -764 119 -744
rect 149 -764 159 -744
rect 90 -776 159 -764
rect 199 -744 269 -734
rect 199 -764 209 -744
rect 239 -764 269 -744
rect 199 -776 269 -764
rect 284 -744 389 -734
rect 284 -764 309 -744
rect 339 -764 389 -744
rect 284 -776 389 -764
rect 404 -744 502 -734
rect 404 -764 429 -744
rect 459 -764 502 -744
rect 404 -776 502 -764
rect 517 -744 612 -734
rect 517 -764 552 -744
rect 582 -764 612 -744
rect 517 -776 612 -764
rect 627 -744 710 -734
rect 627 -764 670 -744
rect 700 -764 710 -744
rect 627 -776 710 -764
rect 750 -744 820 -734
rect 750 -764 760 -744
rect 790 -764 820 -744
rect 750 -776 820 -764
rect 835 -744 940 -734
rect 835 -764 860 -744
rect 890 -764 940 -744
rect 835 -776 940 -764
rect 955 -744 1020 -734
rect 955 -764 980 -744
rect 1010 -764 1020 -744
rect 955 -776 1020 -764
rect 1061 -744 1131 -734
rect 1061 -764 1071 -744
rect 1101 -764 1131 -744
rect 1061 -776 1131 -764
rect 1146 -744 1211 -734
rect 1146 -764 1171 -744
rect 1201 -764 1211 -744
rect 1146 -776 1211 -764
rect 1250 -744 1320 -734
rect 1250 -764 1260 -744
rect 1290 -764 1320 -744
rect 1250 -776 1320 -764
rect 1335 -744 1400 -734
rect 1335 -764 1360 -744
rect 1390 -764 1400 -744
rect 1335 -776 1400 -764
<< pdiff >>
rect 5 -110 75 -70
rect 5 -170 15 -110
rect 55 -170 75 -110
rect 5 -200 75 -170
rect 90 -110 159 -70
rect 90 -170 109 -110
rect 149 -170 159 -110
rect 90 -200 159 -170
rect 199 -110 269 -70
rect 199 -170 209 -110
rect 249 -170 269 -110
rect 199 -200 269 -170
rect 284 -110 389 -70
rect 284 -170 309 -110
rect 349 -170 389 -110
rect 284 -200 389 -170
rect 404 -110 502 -70
rect 404 -170 419 -110
rect 459 -170 502 -110
rect 404 -200 502 -170
rect 517 -110 612 -70
rect 517 -170 542 -110
rect 582 -170 612 -110
rect 517 -200 612 -170
rect 627 -110 710 -70
rect 627 -170 660 -110
rect 700 -170 710 -110
rect 627 -200 710 -170
rect 750 -110 820 -70
rect 750 -170 760 -110
rect 800 -170 820 -110
rect 750 -200 820 -170
rect 835 -110 940 -70
rect 835 -170 850 -110
rect 890 -170 940 -110
rect 835 -200 940 -170
rect 955 -110 1020 -70
rect 955 -170 970 -110
rect 1010 -170 1020 -110
rect 955 -200 1020 -170
rect 1061 -110 1131 -70
rect 1061 -170 1071 -110
rect 1111 -170 1131 -110
rect 1061 -200 1131 -170
rect 1146 -110 1211 -70
rect 1146 -170 1161 -110
rect 1201 -170 1211 -110
rect 1146 -200 1211 -170
rect 1250 -110 1320 -70
rect 1250 -170 1260 -110
rect 1300 -170 1320 -110
rect 1250 -200 1320 -170
rect 1335 -110 1400 -70
rect 1335 -170 1350 -110
rect 1390 -170 1400 -110
rect 1335 -200 1400 -170
<< ndiffc >>
rect 15 -764 45 -744
rect 119 -764 149 -744
rect 209 -764 239 -744
rect 309 -764 339 -744
rect 429 -764 459 -744
rect 552 -764 582 -744
rect 670 -764 700 -744
rect 760 -764 790 -744
rect 860 -764 890 -744
rect 980 -764 1010 -744
rect 1071 -764 1101 -744
rect 1171 -764 1201 -744
rect 1260 -764 1290 -744
rect 1360 -764 1390 -744
<< pdiffc >>
rect 15 -170 55 -110
rect 109 -170 149 -110
rect 209 -170 249 -110
rect 309 -170 349 -110
rect 419 -170 459 -110
rect 542 -170 582 -110
rect 660 -170 700 -110
rect 760 -170 800 -110
rect 850 -170 890 -110
rect 970 -170 1010 -110
rect 1071 -170 1111 -110
rect 1161 -170 1201 -110
rect 1260 -170 1300 -110
rect 1350 -170 1390 -110
<< psubdiff >>
rect -15 -954 55 -934
rect -15 -984 5 -954
rect 35 -984 55 -954
rect -15 -1004 55 -984
rect 85 -954 159 -934
rect 85 -984 109 -954
rect 139 -984 159 -954
rect 85 -1004 159 -984
rect 189 -954 259 -934
rect 189 -984 209 -954
rect 239 -984 259 -954
rect 189 -1004 259 -984
rect 289 -954 379 -934
rect 289 -984 309 -954
rect 339 -984 379 -954
rect 289 -1004 379 -984
rect 409 -954 492 -934
rect 409 -984 429 -954
rect 459 -984 492 -954
rect 409 -1004 492 -984
rect 522 -954 602 -934
rect 522 -984 552 -954
rect 582 -984 602 -954
rect 522 -1004 602 -984
rect 632 -954 710 -934
rect 632 -984 660 -954
rect 690 -984 710 -954
rect 632 -1004 710 -984
rect 740 -954 810 -934
rect 740 -984 760 -954
rect 790 -984 810 -954
rect 740 -1004 810 -984
rect 840 -954 910 -934
rect 840 -984 860 -954
rect 890 -984 910 -954
rect 840 -1004 910 -984
rect 940 -954 1010 -934
rect 940 -984 960 -954
rect 990 -984 1010 -954
rect 940 -1004 1010 -984
rect 1040 -954 1110 -934
rect 1040 -984 1060 -954
rect 1090 -984 1110 -954
rect 1040 -1004 1110 -984
rect 1140 -954 1210 -934
rect 1140 -984 1160 -954
rect 1190 -984 1210 -954
rect 1140 -1004 1210 -984
rect 1240 -954 1310 -934
rect 1240 -984 1260 -954
rect 1290 -984 1310 -954
rect 1240 -1004 1310 -984
rect 1340 -954 1410 -934
rect 1340 -984 1360 -954
rect 1390 -984 1410 -954
rect 1340 -1004 1410 -984
<< nsubdiff >>
rect -15 250 65 270
rect -15 210 5 250
rect 45 210 65 250
rect -15 190 65 210
rect 95 250 179 270
rect 95 210 119 250
rect 159 210 179 250
rect 95 190 179 210
rect 209 250 289 270
rect 209 210 229 250
rect 269 210 289 250
rect 209 190 289 210
rect 319 250 419 270
rect 319 210 339 250
rect 399 210 419 250
rect 319 190 419 210
rect 449 250 552 270
rect 449 210 469 250
rect 522 210 552 250
rect 449 190 552 210
rect 582 250 670 270
rect 582 210 602 250
rect 642 210 670 250
rect 582 190 670 210
rect 700 250 780 270
rect 700 210 720 250
rect 760 210 780 250
rect 700 190 780 210
rect 810 250 890 270
rect 810 210 830 250
rect 870 210 890 250
rect 810 190 890 210
rect 920 250 1000 270
rect 920 210 940 250
rect 980 210 1000 250
rect 920 190 1000 210
rect 1030 250 1110 270
rect 1030 210 1050 250
rect 1090 210 1110 250
rect 1030 190 1110 210
rect 1140 250 1220 270
rect 1140 210 1160 250
rect 1200 210 1220 250
rect 1140 190 1220 210
rect 1250 250 1330 270
rect 1250 210 1270 250
rect 1310 210 1330 250
rect 1250 190 1330 210
rect 1360 250 1440 270
rect 1360 210 1380 250
rect 1420 210 1440 250
rect 1360 190 1440 210
rect -15 140 65 160
rect -15 100 5 140
rect 45 100 65 140
rect -15 80 65 100
rect 95 140 179 160
rect 95 100 119 140
rect 159 100 179 140
rect 95 80 179 100
rect 209 140 289 160
rect 209 100 229 140
rect 269 100 289 140
rect 209 80 289 100
rect 319 140 419 160
rect 319 100 339 140
rect 399 100 419 140
rect 319 80 419 100
rect 449 140 552 160
rect 449 100 469 140
rect 522 100 552 140
rect 449 80 552 100
rect 582 140 670 160
rect 582 100 602 140
rect 642 100 670 140
rect 582 80 670 100
rect 700 140 780 160
rect 700 100 720 140
rect 760 100 780 140
rect 700 80 780 100
rect 810 140 890 160
rect 810 100 830 140
rect 870 100 890 140
rect 810 80 890 100
rect 920 140 1000 160
rect 920 100 940 140
rect 980 100 1000 140
rect 920 80 1000 100
rect 1030 140 1110 160
rect 1030 100 1050 140
rect 1090 100 1110 140
rect 1030 80 1110 100
rect 1140 140 1220 160
rect 1140 100 1160 140
rect 1200 100 1220 140
rect 1140 80 1220 100
rect 1250 140 1330 160
rect 1250 100 1270 140
rect 1310 100 1330 140
rect 1250 80 1330 100
rect 1360 140 1440 160
rect 1360 100 1380 140
rect 1420 100 1440 140
rect 1360 80 1440 100
<< psubdiffcont >>
rect 5 -984 35 -954
rect 109 -984 139 -954
rect 209 -984 239 -954
rect 309 -984 339 -954
rect 429 -984 459 -954
rect 552 -984 582 -954
rect 660 -984 690 -954
rect 760 -984 790 -954
rect 860 -984 890 -954
rect 960 -984 990 -954
rect 1060 -984 1090 -954
rect 1160 -984 1190 -954
rect 1260 -984 1290 -954
rect 1360 -984 1390 -954
<< nsubdiffcont >>
rect 5 210 45 250
rect 119 210 159 250
rect 229 210 269 250
rect 339 210 399 250
rect 469 210 522 250
rect 602 210 642 250
rect 720 210 760 250
rect 830 210 870 250
rect 940 210 980 250
rect 1050 210 1090 250
rect 1160 210 1200 250
rect 1270 210 1310 250
rect 1380 210 1420 250
rect 5 100 45 140
rect 119 100 159 140
rect 229 100 269 140
rect 339 100 399 140
rect 469 100 522 140
rect 602 100 642 140
rect 720 100 760 140
rect 830 100 870 140
rect 940 100 980 140
rect 1050 100 1090 140
rect 1160 100 1200 140
rect 1270 100 1310 140
rect 1380 100 1420 140
<< poly >>
rect 75 -70 90 -50
rect 269 -70 284 -50
rect 389 -70 404 -50
rect 502 -70 517 -50
rect 612 -70 627 -50
rect 820 -70 835 -50
rect 940 -70 955 -50
rect 1131 -70 1146 -50
rect 1320 -70 1335 -50
rect 75 -525 90 -200
rect 269 -480 284 -200
rect 389 -263 404 -200
rect 502 -220 517 -200
rect 612 -220 627 -200
rect 486 -232 627 -220
rect 486 -258 496 -232
rect 522 -240 627 -232
rect 522 -258 531 -240
rect 359 -279 409 -263
rect 486 -270 531 -258
rect 359 -307 370 -279
rect 398 -307 409 -279
rect 359 -313 409 -307
rect 820 -330 835 -200
rect 940 -262 955 -200
rect 910 -278 960 -262
rect 910 -306 921 -278
rect 949 -306 960 -278
rect 910 -312 960 -306
rect 790 -340 835 -330
rect 790 -360 800 -340
rect 820 -360 835 -340
rect 790 -370 835 -360
rect 239 -490 284 -480
rect 239 -510 249 -490
rect 269 -510 284 -490
rect 239 -520 284 -510
rect 47 -537 92 -525
rect 47 -563 57 -537
rect 83 -563 92 -537
rect 47 -575 92 -563
rect 75 -734 90 -575
rect 269 -734 284 -520
rect 367 -541 412 -529
rect 367 -567 377 -541
rect 403 -567 412 -541
rect 367 -579 412 -567
rect 389 -734 404 -579
rect 599 -660 650 -644
rect 599 -688 611 -660
rect 639 -688 650 -660
rect 599 -694 650 -688
rect 502 -714 627 -694
rect 502 -734 517 -714
rect 612 -734 627 -714
rect 820 -734 835 -370
rect 1131 -430 1146 -200
rect 1320 -320 1335 -200
rect 1290 -330 1335 -320
rect 1290 -350 1300 -330
rect 1320 -350 1335 -330
rect 1290 -360 1335 -350
rect 1101 -440 1146 -430
rect 1101 -460 1111 -440
rect 1131 -460 1146 -440
rect 1101 -470 1146 -460
rect 915 -540 960 -528
rect 915 -566 925 -540
rect 951 -566 960 -540
rect 915 -578 960 -566
rect 940 -734 955 -578
rect 1131 -734 1146 -470
rect 1320 -734 1335 -360
rect 75 -794 90 -776
rect 269 -794 284 -776
rect 389 -794 404 -776
rect 502 -794 517 -776
rect 612 -794 627 -776
rect 820 -794 835 -776
rect 940 -794 955 -776
rect 1131 -794 1146 -776
rect 1320 -794 1335 -776
<< polycont >>
rect 496 -258 522 -232
rect 370 -307 398 -279
rect 921 -306 949 -278
rect 800 -360 820 -340
rect 249 -510 269 -490
rect 57 -563 83 -537
rect 377 -567 403 -541
rect 611 -688 639 -660
rect 1300 -350 1320 -330
rect 1111 -460 1131 -440
rect 925 -566 951 -540
<< locali >>
rect -55 250 1458 290
rect -55 210 5 250
rect 45 210 119 250
rect 159 210 229 250
rect 269 210 339 250
rect 399 210 469 250
rect 522 210 602 250
rect 642 210 720 250
rect 760 210 830 250
rect 870 210 940 250
rect 980 210 1050 250
rect 1090 210 1160 250
rect 1200 210 1270 250
rect 1310 210 1380 250
rect 1420 210 1458 250
rect -55 140 1458 210
rect -55 100 5 140
rect 45 100 119 140
rect 159 100 229 140
rect 269 100 339 140
rect 399 100 469 140
rect 522 100 602 140
rect 642 100 720 140
rect 760 100 830 140
rect 870 100 940 140
rect 980 100 1050 140
rect 1090 100 1160 140
rect 1200 100 1270 140
rect 1310 100 1380 140
rect 1420 100 1458 140
rect -55 60 1458 100
rect 15 -70 45 60
rect 209 -70 239 60
rect 760 -70 790 60
rect 1071 -70 1101 60
rect 1260 -70 1290 60
rect 5 -110 55 -70
rect 5 -170 15 -110
rect 5 -200 55 -170
rect 109 -110 159 -70
rect 149 -170 159 -110
rect 109 -200 159 -170
rect 199 -110 249 -70
rect 199 -170 209 -110
rect 199 -200 249 -170
rect 299 -110 349 -70
rect 299 -170 309 -110
rect 299 -200 349 -170
rect 419 -110 469 -70
rect 459 -170 469 -110
rect 419 -200 469 -170
rect 542 -110 592 -70
rect 582 -170 592 -110
rect 542 -200 592 -170
rect 660 -110 710 -70
rect 700 -170 710 -110
rect 660 -200 710 -170
rect 750 -110 800 -70
rect 750 -170 760 -110
rect 750 -200 800 -170
rect 850 -110 900 -70
rect 890 -170 900 -110
rect 850 -200 900 -170
rect 970 -110 1020 -70
rect 1010 -170 1020 -110
rect 970 -200 1020 -170
rect 1061 -110 1111 -70
rect 1061 -170 1071 -110
rect 1061 -200 1111 -170
rect 1161 -110 1211 -70
rect 1201 -170 1211 -110
rect 1161 -200 1211 -170
rect 1250 -110 1300 -70
rect 1250 -170 1260 -110
rect 1250 -200 1300 -170
rect 1350 -110 1400 -70
rect 1390 -170 1400 -110
rect 1350 -200 1400 -170
rect 119 -380 149 -200
rect 309 -330 339 -200
rect 359 -279 409 -263
rect 359 -307 370 -279
rect 398 -307 409 -279
rect 359 -313 409 -307
rect 309 -340 349 -330
rect 309 -360 319 -340
rect 339 -360 349 -340
rect 309 -370 349 -360
rect 114 -391 164 -380
rect 114 -419 125 -391
rect 153 -419 164 -391
rect 114 -430 164 -419
rect 47 -537 92 -525
rect 47 -547 57 -537
rect 16 -563 57 -547
rect 83 -563 92 -537
rect 16 -572 92 -563
rect 47 -575 92 -572
rect 119 -734 149 -430
rect 239 -490 284 -480
rect 239 -510 249 -490
rect 269 -510 284 -490
rect 239 -520 284 -510
rect 309 -734 339 -370
rect 429 -430 459 -200
rect 486 -232 531 -220
rect 486 -258 496 -232
rect 522 -258 531 -232
rect 486 -270 531 -258
rect 429 -440 469 -430
rect 429 -460 439 -440
rect 459 -460 469 -440
rect 429 -470 469 -460
rect 367 -541 412 -529
rect 367 -567 377 -541
rect 403 -567 412 -541
rect 367 -579 412 -567
rect 429 -734 459 -470
rect 552 -580 582 -200
rect 670 -480 700 -200
rect 790 -340 835 -330
rect 790 -360 800 -340
rect 820 -360 835 -340
rect 790 -370 835 -360
rect 670 -490 710 -480
rect 670 -510 680 -490
rect 700 -510 710 -490
rect 670 -520 710 -510
rect 552 -590 592 -580
rect 552 -610 562 -590
rect 582 -610 592 -590
rect 552 -620 592 -610
rect 552 -734 582 -620
rect 599 -660 650 -644
rect 599 -688 611 -660
rect 639 -688 650 -660
rect 599 -694 650 -688
rect 670 -734 700 -520
rect 860 -734 890 -200
rect 910 -278 960 -262
rect 910 -306 921 -278
rect 949 -306 960 -278
rect 910 -312 960 -306
rect 980 -480 1010 -200
rect 1171 -320 1201 -200
rect 1171 -330 1211 -320
rect 1290 -330 1335 -320
rect 1171 -350 1181 -330
rect 1201 -350 1300 -330
rect 1320 -350 1335 -330
rect 1171 -360 1335 -350
rect 1101 -440 1146 -430
rect 1101 -460 1111 -440
rect 1131 -460 1146 -440
rect 1101 -470 1146 -460
rect 980 -490 1020 -480
rect 980 -510 990 -490
rect 1010 -510 1020 -490
rect 980 -520 1020 -510
rect 915 -540 960 -528
rect 915 -566 925 -540
rect 951 -566 960 -540
rect 915 -578 960 -566
rect 980 -734 1010 -520
rect 1171 -734 1201 -360
rect 1360 -581 1390 -200
rect 1360 -591 1400 -581
rect 1360 -611 1370 -591
rect 1390 -611 1400 -591
rect 1360 -621 1400 -611
rect 1360 -734 1390 -621
rect 5 -744 55 -734
rect 5 -764 15 -744
rect 45 -764 55 -744
rect 5 -776 55 -764
rect 109 -744 159 -734
rect 109 -764 119 -744
rect 149 -764 159 -744
rect 109 -776 159 -764
rect 199 -744 249 -734
rect 199 -764 209 -744
rect 239 -764 249 -744
rect 199 -776 249 -764
rect 299 -744 349 -734
rect 299 -764 309 -744
rect 339 -764 349 -744
rect 299 -776 349 -764
rect 419 -744 469 -734
rect 419 -764 429 -744
rect 459 -764 469 -744
rect 419 -776 469 -764
rect 542 -744 592 -734
rect 542 -764 552 -744
rect 582 -764 592 -744
rect 542 -776 592 -764
rect 660 -744 710 -734
rect 660 -764 670 -744
rect 700 -764 710 -744
rect 660 -776 710 -764
rect 750 -744 800 -734
rect 750 -764 760 -744
rect 790 -764 800 -744
rect 750 -776 800 -764
rect 850 -744 900 -734
rect 850 -764 860 -744
rect 890 -764 900 -744
rect 850 -776 900 -764
rect 970 -744 1020 -734
rect 970 -764 980 -744
rect 1010 -764 1020 -744
rect 970 -776 1020 -764
rect 1061 -744 1111 -734
rect 1061 -764 1071 -744
rect 1101 -764 1111 -744
rect 1061 -776 1111 -764
rect 1161 -744 1211 -734
rect 1161 -764 1171 -744
rect 1201 -764 1211 -744
rect 1161 -776 1211 -764
rect 1250 -744 1300 -734
rect 1250 -764 1260 -744
rect 1290 -764 1300 -744
rect 1250 -776 1300 -764
rect 1350 -744 1400 -734
rect 1350 -764 1360 -744
rect 1390 -764 1400 -744
rect 1350 -776 1400 -764
rect 15 -914 45 -776
rect 209 -914 239 -776
rect 760 -914 790 -776
rect 1071 -914 1101 -776
rect 1260 -914 1290 -776
rect -55 -954 1480 -914
rect -55 -984 5 -954
rect 35 -984 109 -954
rect 139 -984 209 -954
rect 239 -984 309 -954
rect 339 -984 429 -954
rect 459 -984 552 -954
rect 582 -984 660 -954
rect 690 -984 760 -954
rect 790 -984 860 -954
rect 890 -984 960 -954
rect 990 -984 1060 -954
rect 1090 -984 1160 -954
rect 1190 -984 1260 -954
rect 1290 -984 1360 -954
rect 1390 -984 1480 -954
rect -55 -1034 1480 -984
<< viali >>
rect 370 -307 398 -279
rect 319 -360 339 -340
rect 125 -419 153 -391
rect 57 -563 83 -537
rect 249 -510 269 -490
rect 496 -258 522 -232
rect 439 -460 459 -440
rect 377 -567 403 -541
rect 800 -360 820 -340
rect 680 -510 700 -490
rect 562 -610 582 -590
rect 611 -688 639 -660
rect 921 -306 949 -278
rect 1181 -350 1201 -330
rect 1300 -350 1320 -330
rect 1111 -460 1131 -440
rect 990 -510 1010 -490
rect 925 -566 951 -540
rect 1370 -611 1390 -591
<< metal1 >>
rect 486 -232 531 -220
rect 486 -258 496 -232
rect 522 -258 531 -232
rect 359 -279 409 -263
rect 486 -270 531 -258
rect 359 -307 370 -279
rect 398 -307 409 -279
rect 359 -313 409 -307
rect 910 -278 960 -262
rect 910 -306 921 -278
rect 949 -306 960 -278
rect 910 -312 960 -306
rect 1171 -330 1211 -320
rect 309 -340 349 -330
rect 790 -340 835 -330
rect 309 -360 319 -340
rect 339 -360 800 -340
rect 820 -360 835 -340
rect 1171 -350 1181 -330
rect 1201 -350 1211 -330
rect 1171 -360 1211 -350
rect 1290 -330 1335 -320
rect 1290 -350 1300 -330
rect 1320 -350 1458 -330
rect 1290 -360 1458 -350
rect 309 -370 835 -360
rect 114 -391 164 -380
rect 114 -419 125 -391
rect 153 -419 164 -391
rect 114 -430 164 -419
rect 429 -440 1146 -430
rect 429 -460 439 -440
rect 459 -460 1111 -440
rect 1131 -460 1146 -440
rect 429 -470 469 -460
rect 1101 -470 1146 -460
rect 239 -484 284 -480
rect 670 -484 710 -480
rect 980 -484 1020 -480
rect 239 -490 1020 -484
rect 239 -510 249 -490
rect 269 -510 680 -490
rect 700 -510 990 -490
rect 1010 -510 1020 -490
rect 239 -514 1020 -510
rect 239 -520 284 -514
rect 670 -520 710 -514
rect 980 -520 1020 -514
rect 47 -537 92 -525
rect 47 -563 57 -537
rect 83 -563 92 -537
rect 47 -575 92 -563
rect 367 -541 412 -529
rect 367 -567 377 -541
rect 403 -567 412 -541
rect 367 -579 412 -567
rect 915 -540 960 -528
rect 915 -566 925 -540
rect 951 -566 960 -540
rect 915 -578 960 -566
rect 552 -590 592 -580
rect 552 -610 562 -590
rect 582 -595 592 -590
rect 1360 -591 1400 -581
rect 1360 -595 1370 -591
rect 582 -610 1370 -595
rect 552 -611 1370 -610
rect 1390 -611 1400 -591
rect 552 -620 1400 -611
rect 1360 -621 1400 -620
rect 599 -660 650 -644
rect 599 -688 611 -660
rect 639 -688 650 -660
rect 599 -694 650 -688
<< via1 >>
rect 496 -258 522 -232
rect 370 -307 398 -279
rect 921 -306 949 -278
rect 125 -419 153 -391
rect 57 -563 83 -537
rect 377 -567 403 -541
rect 925 -566 951 -540
rect 611 -688 639 -660
<< metal2 >>
rect 486 -232 531 -220
rect 486 -258 496 -232
rect 522 -258 531 -232
rect 359 -279 409 -263
rect 486 -270 531 -258
rect 359 -307 370 -279
rect 398 -307 409 -279
rect 359 -313 409 -307
rect 114 -391 164 -380
rect 114 -419 125 -391
rect 153 -419 164 -391
rect 114 -430 164 -419
rect 47 -537 92 -525
rect 47 -563 57 -537
rect 83 -540 92 -537
rect 367 -540 412 -529
rect 500 -540 530 -270
rect 910 -278 960 -262
rect 910 -306 921 -278
rect 949 -306 960 -278
rect 910 -312 960 -306
rect 915 -540 960 -528
rect 83 -541 925 -540
rect 83 -563 377 -541
rect 47 -567 377 -563
rect 403 -566 925 -541
rect 951 -566 960 -540
rect 403 -567 960 -566
rect 47 -570 960 -567
rect 47 -575 92 -570
rect 367 -579 412 -570
rect 915 -578 960 -570
rect 599 -660 650 -644
rect 599 -688 611 -660
rect 639 -688 650 -660
rect 599 -694 650 -688
<< via2 >>
rect 370 -307 398 -279
rect 125 -419 153 -391
rect 921 -306 949 -278
rect 611 -688 639 -660
<< metal3 >>
rect 359 -279 409 -263
rect 910 -270 960 -262
rect 359 -307 370 -279
rect 398 -307 409 -279
rect 359 -313 409 -307
rect 369 -380 409 -313
rect 610 -278 960 -270
rect 610 -306 921 -278
rect 949 -306 960 -278
rect 610 -310 960 -306
rect 610 -380 650 -310
rect 910 -312 960 -310
rect 114 -391 650 -380
rect 114 -419 125 -391
rect 153 -419 650 -391
rect 114 -420 650 -419
rect 114 -430 164 -420
rect 610 -644 650 -420
rect 599 -660 650 -644
rect 599 -688 611 -660
rect 639 -688 650 -660
rect 599 -694 650 -688
<< labels >>
rlabel locali 709 -1027 757 -1008 1 gnd!
rlabel locali 673 164 693 176 1 vdd
rlabel locali 22 -567 35 -559 1 clk
rlabel metal1 1415 -358 1453 -338 1 q
<< end >>
