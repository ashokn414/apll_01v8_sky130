***pfd circuit***
.param L=0.15
.param W=0.42
.include "/home/ashok/sky130_fd_pr/models/corners/tt.spice"
.include "/home/ashok/Desktop/tools/spice_exp/ashvsdpll/inverter.lib"
.include "/home/ashok/Desktop/tools/spice_exp/ashvsdpll/nand1.lib"
.include "/home/ashok/Desktop/tools/spice_exp/ashvsdpll/nand2.lib"
.include "/home/ashok/Desktop/tools/spice_exp/ashvsdpll/nand3.lib"

XX1 N001 N005 N002 vddd 0 nand1
XX2 N002 N008 N006 vddd 0 nand1
XX3 N006 N007 N008 vddd 0 nand1
XX4 N007 N010 N011 vddd 0 nand1
XX5 N011 N009 N010 vddd 0 nand1
XX6 N013 N012 N009 vddd 0 nand1
XX7 f_clk_in N005 vddd 0 inverter
XX8 f_VCO N013 vddd 0 inverter
XX9 N002 N003 vddd 0 inverter
XX10 N003 N004 vddd 0 inverter
XX11 N009 N014 vddd 0 inverter
XX12 N014 N015 vddd 0 inverter
XX13 N004 N006 N007 N001 vddd 0 nand2
XX14 N007 N010 N015 N012 vddd 0 nand2
XX15 N012 down vddd 0 inverter
XX16 N006 N002 N009 N010 vddd 0 N007 nand3
XX17 N001 up vddd 0 inverter
V3 vddd 0 1.8

***set supply ***

Vin1 f_clk_in 0 0 pulse(0 1 0 100p 100p 5n 10n) 
Vin2 f_VCO 0 0 pulse(0 1 2n 100p 100p 5n 9n)
 
.op
.tran 10p 50n
.end
