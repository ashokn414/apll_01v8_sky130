magic
tech sky130A
timestamp 1605793028
<< nwell >>
rect 2010 4041 2530 4220
rect 1690 4040 2530 4041
rect 1550 3600 2530 4040
rect 1690 3599 2530 3600
<< nmos >>
rect 1810 4236 1825 4278
rect 1890 4236 1905 4278
rect 1810 3362 1825 3404
rect 1890 3362 1905 3404
rect 2070 3375 2112 3390
rect 2290 3355 2332 3370
rect 2000 2996 2015 3220
rect 2165 3178 2180 3220
<< pmos >>
rect 2100 4139 2184 4154
rect 2256 4053 2340 4068
rect 1810 3929 1825 4013
rect 1890 3929 1905 4013
rect 1810 3627 1825 3711
rect 1890 3627 1905 3711
rect 2120 3625 2135 4025
rect 2200 3625 2215 3709
<< ndiff >>
rect 1760 4270 1810 4278
rect 1760 4246 1768 4270
rect 1792 4246 1810 4270
rect 1760 4236 1810 4246
rect 1825 4270 1890 4278
rect 1825 4246 1848 4270
rect 1872 4246 1890 4270
rect 1825 4236 1890 4246
rect 1905 4270 1960 4278
rect 1905 4246 1928 4270
rect 1952 4246 1960 4270
rect 1905 4236 1960 4246
rect 1759 3404 1800 3405
rect 2070 3432 2112 3440
rect 2070 3408 2078 3432
rect 2102 3408 2112 3432
rect 1759 3396 1810 3404
rect 1759 3370 1766 3396
rect 1792 3370 1810 3396
rect 1759 3362 1810 3370
rect 1825 3394 1890 3404
rect 1825 3370 1848 3394
rect 1872 3370 1890 3394
rect 1825 3362 1890 3370
rect 1905 3394 1960 3404
rect 1905 3370 1928 3394
rect 1952 3370 1960 3394
rect 1905 3362 1960 3370
rect 2070 3390 2112 3408
rect 2289 3414 2333 3422
rect 2289 3388 2298 3414
rect 2324 3388 2333 3414
rect 2289 3380 2333 3388
rect 2070 3352 2112 3375
rect 2290 3370 2332 3380
rect 2070 3328 2078 3352
rect 2102 3328 2112 3352
rect 2070 3320 2112 3328
rect 1945 3220 1986 3221
rect 2290 3340 2332 3355
rect 2289 3332 2332 3340
rect 2289 3300 2298 3332
rect 2324 3300 2332 3332
rect 2289 3290 2332 3300
rect 1945 3212 2000 3220
rect 1945 3030 1952 3212
rect 1978 3030 2000 3212
rect 1945 2996 2000 3030
rect 2015 3211 2165 3220
rect 2015 3029 2077 3211
rect 2103 3178 2165 3211
rect 2180 3210 2255 3220
rect 2180 3186 2223 3210
rect 2247 3186 2255 3210
rect 2180 3178 2255 3186
rect 2103 3029 2110 3178
rect 2015 2996 2110 3029
<< pdiff >>
rect 2100 4196 2184 4202
rect 2100 4176 2123 4196
rect 2158 4176 2184 4196
rect 2100 4154 2184 4176
rect 2100 4118 2184 4139
rect 2100 4098 2123 4118
rect 2158 4098 2184 4118
rect 2100 4088 2184 4098
rect 2256 4114 2340 4118
rect 2256 4085 2276 4114
rect 2316 4085 2340 4114
rect 2256 4068 2340 4085
rect 1760 3987 1810 4013
rect 1760 3954 1766 3987
rect 1793 3954 1810 3987
rect 1760 3929 1810 3954
rect 1825 3989 1890 4013
rect 1825 3949 1843 3989
rect 1873 3949 1890 3989
rect 1825 3929 1890 3949
rect 1905 3989 1960 4013
rect 1905 3949 1923 3989
rect 1953 3949 1960 3989
rect 1905 3929 1960 3949
rect 2070 3987 2120 4025
rect 1760 3685 1810 3711
rect 1760 3652 1766 3685
rect 1793 3652 1810 3685
rect 1760 3627 1810 3652
rect 1825 3691 1890 3711
rect 1825 3651 1843 3691
rect 1873 3651 1890 3691
rect 1825 3627 1890 3651
rect 1905 3687 1960 3711
rect 1905 3647 1923 3687
rect 1953 3647 1960 3687
rect 1905 3627 1960 3647
rect 2070 3650 2076 3987
rect 2103 3650 2120 3987
rect 2070 3625 2120 3650
rect 2135 3984 2190 4025
rect 2135 3647 2156 3984
rect 2183 3709 2190 3984
rect 2256 4031 2340 4053
rect 2256 4005 2281 4031
rect 2316 4005 2340 4031
rect 2256 3998 2340 4005
rect 2183 3647 2200 3709
rect 2135 3625 2200 3647
rect 2215 3685 2270 3709
rect 2215 3645 2233 3685
rect 2263 3645 2270 3685
rect 2215 3625 2270 3645
<< ndiffc >>
rect 1768 4246 1792 4270
rect 1848 4246 1872 4270
rect 1928 4246 1952 4270
rect 2078 3408 2102 3432
rect 1766 3370 1792 3396
rect 1848 3370 1872 3394
rect 1928 3370 1952 3394
rect 2298 3388 2324 3414
rect 2078 3328 2102 3352
rect 2298 3300 2324 3332
rect 1952 3030 1978 3212
rect 2077 3029 2103 3211
rect 2223 3186 2247 3210
<< pdiffc >>
rect 2123 4176 2158 4196
rect 2123 4098 2158 4118
rect 2276 4085 2316 4114
rect 1766 3954 1793 3987
rect 1843 3949 1873 3989
rect 1923 3949 1953 3989
rect 1766 3652 1793 3685
rect 1843 3651 1873 3691
rect 1923 3647 1953 3687
rect 2076 3650 2103 3987
rect 2156 3647 2183 3984
rect 2281 4005 2316 4031
rect 2233 3645 2263 3685
<< psubdiff >>
rect 1488 4387 1850 4397
rect 1488 4347 1510 4387
rect 1550 4347 1580 4387
rect 1620 4347 1650 4387
rect 1690 4347 1720 4387
rect 1760 4347 1790 4387
rect 1830 4347 1850 4387
rect 1930 4387 2330 4397
rect 1488 4337 1850 4347
rect 1930 4347 1950 4387
rect 1990 4347 2020 4387
rect 2060 4347 2090 4387
rect 2130 4347 2160 4387
rect 2200 4347 2230 4387
rect 2270 4347 2330 4387
rect 1930 4337 2330 4347
<< nsubdiff >>
rect 1720 3870 1860 3880
rect 1720 3830 1740 3870
rect 1780 3830 1800 3870
rect 1840 3830 1860 3870
rect 1720 3810 1860 3830
rect 1720 3770 1740 3810
rect 1780 3770 1800 3810
rect 1840 3770 1860 3810
rect 1720 3760 1860 3770
rect 2390 4021 2452 4030
rect 2390 3987 2404 4021
rect 2437 3987 2452 4021
rect 2390 3980 2452 3987
<< psubdiffcont >>
rect 1510 4347 1550 4387
rect 1580 4347 1620 4387
rect 1650 4347 1690 4387
rect 1720 4347 1760 4387
rect 1790 4347 1830 4387
rect 1950 4347 1990 4387
rect 2020 4347 2060 4387
rect 2090 4347 2130 4387
rect 2160 4347 2200 4387
rect 2230 4347 2270 4387
<< nsubdiffcont >>
rect 1740 3830 1780 3870
rect 1800 3830 1840 3870
rect 1740 3770 1780 3810
rect 1800 3770 1840 3810
rect 2404 3987 2437 4021
<< poly >>
rect 1870 4358 1910 4368
rect 1870 4338 1880 4358
rect 1900 4338 1910 4358
rect 1870 4328 1910 4338
rect 1810 4278 1825 4298
rect 1890 4278 1905 4328
rect 1810 4160 1825 4236
rect 1890 4216 1905 4236
rect 1785 4150 1825 4160
rect 1785 4130 1795 4150
rect 1815 4130 1825 4150
rect 1785 4120 1825 4130
rect 2019 4158 2059 4168
rect 2019 4138 2029 4158
rect 2049 4154 2059 4158
rect 2320 4180 2376 4190
rect 2320 4160 2330 4180
rect 2350 4160 2376 4180
rect 2049 4139 2100 4154
rect 2184 4139 2204 4154
rect 2320 4150 2376 4160
rect 2049 4138 2059 4139
rect 2019 4128 2059 4138
rect 1810 4013 1825 4120
rect 2010 4065 2050 4070
rect 2360 4068 2376 4150
rect 2010 4060 2135 4065
rect 2010 4040 2020 4060
rect 2040 4050 2135 4060
rect 2040 4040 2050 4050
rect 1890 4013 1905 4033
rect 2010 4030 2050 4040
rect 2120 4025 2135 4050
rect 2200 4053 2256 4068
rect 2340 4053 2376 4068
rect 1810 3909 1825 3929
rect 1890 3831 1905 3929
rect 1879 3823 1921 3831
rect 1879 3797 1887 3823
rect 1913 3797 1921 3823
rect 1879 3789 1921 3797
rect 1810 3711 1825 3731
rect 1890 3711 1905 3789
rect 1810 3520 1825 3627
rect 1890 3607 1905 3627
rect 2200 3709 2215 4053
rect 2120 3605 2135 3625
rect 2200 3605 2215 3625
rect 1785 3510 1825 3520
rect 1785 3490 1795 3510
rect 1815 3490 1825 3510
rect 1785 3480 1825 3490
rect 1810 3404 1825 3480
rect 2356 3456 2400 3466
rect 1890 3404 1905 3424
rect 2356 3430 2366 3456
rect 2392 3430 2400 3456
rect 1990 3390 2030 3400
rect 2356 3420 2400 3430
rect 1990 3370 2000 3390
rect 2020 3375 2070 3390
rect 2112 3375 2132 3390
rect 2020 3370 2030 3375
rect 1810 3342 1825 3362
rect 1890 3332 1905 3362
rect 1990 3360 2030 3370
rect 2370 3370 2385 3420
rect 1880 3324 1922 3332
rect 1880 3298 1888 3324
rect 1914 3298 1922 3324
rect 2165 3355 2290 3370
rect 2332 3355 2385 3370
rect 1880 3290 1922 3298
rect 1990 3274 2032 3280
rect 1990 3251 1999 3274
rect 2021 3251 2032 3274
rect 1990 3242 2032 3251
rect 2000 3220 2015 3242
rect 2165 3220 2180 3355
rect 2165 3158 2180 3178
rect 2000 2975 2015 2996
<< polycont >>
rect 1880 4338 1900 4358
rect 1795 4130 1815 4150
rect 2029 4138 2049 4158
rect 2330 4160 2350 4180
rect 2020 4040 2040 4060
rect 1887 3797 1913 3823
rect 1795 3490 1815 3510
rect 2366 3430 2392 3456
rect 2000 3370 2020 3390
rect 1888 3298 1914 3324
rect 1999 3251 2021 3274
<< locali >>
rect 1420 4407 1517 4408
rect 1420 4387 2340 4407
rect 1420 4347 1510 4387
rect 1550 4347 1580 4387
rect 1620 4347 1650 4387
rect 1690 4347 1720 4387
rect 1760 4347 1790 4387
rect 1830 4358 1950 4387
rect 1830 4347 1880 4358
rect 1420 4338 1880 4347
rect 1900 4347 1950 4358
rect 1990 4347 2020 4387
rect 2060 4347 2090 4387
rect 2130 4347 2160 4387
rect 2200 4347 2230 4387
rect 2270 4347 2340 4387
rect 1900 4338 2340 4347
rect 1420 4328 2340 4338
rect 1420 3390 1460 4328
rect 1760 4278 1790 4328
rect 1760 4270 1800 4278
rect 1760 4246 1768 4270
rect 1792 4246 1800 4270
rect 1760 4236 1800 4246
rect 1840 4270 1880 4278
rect 1840 4246 1848 4270
rect 1872 4246 1880 4270
rect 1840 4236 1880 4246
rect 1920 4270 1960 4278
rect 1920 4246 1928 4270
rect 1952 4246 1960 4270
rect 1920 4236 1960 4246
rect 1785 4150 1825 4160
rect 1785 4130 1795 4150
rect 1815 4130 1825 4150
rect 1785 4120 1825 4130
rect 1850 4013 1880 4236
rect 1930 4013 1960 4236
rect 2100 4196 2184 4202
rect 2100 4176 2123 4196
rect 2158 4176 2184 4196
rect 2100 4168 2184 4176
rect 2290 4190 2340 4328
rect 2290 4180 2360 4190
rect 2019 4158 2059 4168
rect 2019 4138 2029 4158
rect 2049 4138 2059 4158
rect 2019 4128 2059 4138
rect 2290 4160 2330 4180
rect 2350 4160 2360 4180
rect 2290 4150 2360 4160
rect 2100 4118 2184 4128
rect 2290 4118 2340 4150
rect 2100 4098 2123 4118
rect 2158 4098 2184 4118
rect 2100 4088 2184 4098
rect 2256 4114 2340 4118
rect 2256 4085 2276 4114
rect 2316 4085 2340 4114
rect 2256 4078 2340 4085
rect 1760 3987 1800 4013
rect 1760 3954 1766 3987
rect 1793 3954 1800 3987
rect 1760 3929 1800 3954
rect 1840 3989 1880 4013
rect 1840 3949 1843 3989
rect 1873 3949 1880 3989
rect 1840 3929 1880 3949
rect 1920 3989 1960 4013
rect 1920 3949 1923 3989
rect 1953 3970 1960 3989
rect 2010 4060 2050 4070
rect 2010 4040 2020 4060
rect 2040 4040 2050 4060
rect 2010 4030 2050 4040
rect 2256 4031 2520 4038
rect 2010 3970 2040 4030
rect 1953 3949 2040 3970
rect 1920 3940 2040 3949
rect 2070 3987 2110 4025
rect 1920 3929 1960 3940
rect 1760 3890 1790 3929
rect 1589 3870 1950 3890
rect 1589 3853 1740 3870
rect 1589 3827 1627 3853
rect 1653 3830 1740 3853
rect 1780 3830 1800 3870
rect 1840 3830 1950 3870
rect 1653 3827 1950 3830
rect 1589 3823 1950 3827
rect 1589 3810 1887 3823
rect 1589 3770 1740 3810
rect 1780 3770 1800 3810
rect 1840 3797 1887 3810
rect 1913 3797 1950 3823
rect 1840 3770 1950 3797
rect 1589 3750 1950 3770
rect 1760 3711 1790 3750
rect 1760 3685 1800 3711
rect 1760 3652 1766 3685
rect 1793 3652 1800 3685
rect 1760 3627 1800 3652
rect 1840 3691 1880 3711
rect 1840 3651 1843 3691
rect 1873 3651 1880 3691
rect 1840 3627 1880 3651
rect 1920 3687 1960 3711
rect 1920 3647 1923 3687
rect 1953 3647 1960 3687
rect 1920 3627 1960 3647
rect 1785 3510 1825 3520
rect 1785 3490 1795 3510
rect 1815 3490 1825 3510
rect 1785 3480 1825 3490
rect 1580 3399 1630 3410
rect 1580 3390 1592 3399
rect 1420 3372 1592 3390
rect 1618 3372 1630 3399
rect 1420 3360 1630 3372
rect 1759 3396 1800 3405
rect 1850 3404 1880 3627
rect 1930 3404 1960 3627
rect 2070 3650 2076 3987
rect 2103 3650 2110 3987
rect 2070 3625 2110 3650
rect 2150 3984 2190 4025
rect 2256 4005 2281 4031
rect 2316 4022 2520 4031
rect 2316 4021 2467 4022
rect 2316 4005 2404 4021
rect 2256 3998 2404 4005
rect 2340 3997 2404 3998
rect 2150 3647 2156 3984
rect 2183 3647 2190 3984
rect 2390 3987 2404 3997
rect 2437 3996 2467 4021
rect 2493 3996 2520 4022
rect 2437 3987 2520 3996
rect 2390 3970 2520 3987
rect 2150 3625 2190 3647
rect 2230 3685 2270 3709
rect 2230 3645 2233 3685
rect 2263 3655 2270 3685
rect 2263 3645 2450 3655
rect 2230 3625 2450 3645
rect 2356 3456 2400 3466
rect 1759 3370 1766 3396
rect 1792 3370 1800 3396
rect 1759 3362 1800 3370
rect 1840 3394 1880 3404
rect 1840 3370 1848 3394
rect 1872 3370 1880 3394
rect 1840 3362 1880 3370
rect 1920 3394 1960 3404
rect 2070 3432 2112 3440
rect 2070 3408 2078 3432
rect 2102 3408 2112 3432
rect 2356 3430 2366 3456
rect 2392 3430 2400 3456
rect 2070 3400 2112 3408
rect 2289 3414 2333 3422
rect 2356 3420 2400 3430
rect 1920 3370 1928 3394
rect 1952 3370 1960 3394
rect 1920 3362 1960 3370
rect 1990 3390 2030 3400
rect 1990 3370 2000 3390
rect 2020 3370 2030 3390
rect 2289 3388 2298 3414
rect 2324 3388 2333 3414
rect 2289 3380 2333 3388
rect 1990 3360 2030 3370
rect 2070 3352 2112 3360
rect 1880 3324 1922 3332
rect 1880 3298 1888 3324
rect 1914 3298 1922 3324
rect 2070 3328 2078 3352
rect 2102 3328 2112 3352
rect 2070 3320 2112 3328
rect 2289 3332 2332 3340
rect 1880 3290 1922 3298
rect 2289 3300 2298 3332
rect 2324 3300 2332 3332
rect 2289 3290 2332 3300
rect 1990 3274 2032 3280
rect 1990 3251 1999 3274
rect 2021 3251 2032 3274
rect 1990 3242 2032 3251
rect 1945 3212 1986 3221
rect 1945 3030 1952 3212
rect 1978 3030 1986 3212
rect 1945 2996 1986 3030
rect 2070 3211 2110 3220
rect 2070 3029 2077 3211
rect 2103 3029 2110 3211
rect 2215 3210 2255 3220
rect 2215 3186 2223 3210
rect 2247 3208 2255 3210
rect 2420 3208 2450 3625
rect 2247 3186 2450 3208
rect 2215 3178 2450 3186
rect 2070 2996 2110 3029
<< viali >>
rect 1795 4130 1815 4150
rect 2123 4176 2158 4196
rect 2029 4138 2049 4158
rect 2123 4098 2158 4118
rect 1766 3954 1793 3987
rect 1627 3827 1653 3853
rect 1887 3797 1913 3823
rect 1766 3652 1793 3685
rect 1795 3490 1815 3510
rect 1592 3372 1618 3399
rect 2076 3650 2103 3987
rect 2281 4005 2316 4031
rect 2156 3647 2183 3984
rect 2467 3996 2493 4022
rect 1766 3370 1792 3396
rect 2078 3408 2102 3432
rect 2366 3430 2392 3456
rect 2000 3370 2020 3390
rect 2298 3388 2324 3414
rect 1888 3298 1914 3324
rect 2078 3328 2102 3352
rect 2298 3300 2324 3332
rect 1999 3251 2021 3274
rect 1952 3030 1978 3212
rect 2077 3029 2103 3211
<< metal1 >>
rect 2100 4196 2184 4202
rect 2100 4176 2123 4196
rect 2158 4176 2184 4196
rect 2019 4160 2059 4168
rect 1663 4158 2059 4160
rect 1663 4150 2029 4158
rect 1663 4130 1795 4150
rect 1815 4138 2029 4150
rect 2049 4138 2059 4158
rect 1815 4130 2059 4138
rect 1785 4120 1825 4130
rect 2019 4128 2059 4130
rect 2100 4118 2184 4176
rect 2100 4098 2123 4118
rect 2158 4098 2184 4118
rect 2100 4088 2184 4098
rect 2150 4025 2180 4088
rect 2256 4031 2340 4038
rect 1760 3987 1800 4013
rect 1760 3954 1766 3987
rect 1793 3954 1800 3987
rect 1760 3929 1800 3954
rect 2070 3987 2110 4025
rect 1620 3853 1660 3860
rect 1620 3827 1627 3853
rect 1653 3827 1660 3853
rect 1620 3820 1660 3827
rect 1879 3823 1921 3831
rect 1879 3797 1887 3823
rect 1913 3797 1921 3823
rect 1879 3789 1921 3797
rect 1760 3685 1800 3711
rect 1760 3652 1766 3685
rect 1793 3652 1800 3685
rect 1760 3627 1800 3652
rect 2070 3650 2076 3987
rect 2103 3650 2110 3987
rect 2070 3625 2110 3650
rect 2150 3984 2190 4025
rect 2256 4005 2281 4031
rect 2316 4005 2340 4031
rect 2256 3998 2340 4005
rect 2460 4022 2500 4030
rect 2460 3996 2467 4022
rect 2493 3996 2500 4022
rect 2460 3990 2500 3996
rect 2150 3647 2156 3984
rect 2183 3647 2190 3984
rect 2150 3625 2190 3647
rect 1785 3510 1825 3520
rect 1625 3490 1795 3510
rect 1815 3490 2020 3510
rect 1625 3480 2020 3490
rect 1580 3399 1630 3410
rect 1580 3372 1592 3399
rect 1618 3372 1630 3399
rect 1580 3360 1630 3372
rect 1759 3396 1800 3405
rect 1759 3370 1766 3396
rect 1792 3370 1800 3396
rect 1759 3362 1800 3370
rect 1990 3400 2020 3480
rect 2356 3456 2400 3466
rect 2070 3432 2112 3440
rect 2070 3408 2078 3432
rect 2102 3408 2112 3432
rect 2356 3430 2366 3456
rect 2392 3430 2400 3456
rect 2070 3400 2112 3408
rect 2289 3414 2333 3422
rect 2356 3420 2400 3430
rect 1990 3390 2030 3400
rect 1990 3370 2000 3390
rect 2020 3370 2030 3390
rect 1990 3360 2030 3370
rect 2081 3360 2110 3400
rect 2289 3388 2298 3414
rect 2324 3388 2333 3414
rect 2289 3380 2333 3388
rect 1880 3324 1922 3332
rect 1880 3298 1888 3324
rect 1914 3298 1922 3324
rect 1880 3290 1922 3298
rect 1990 3280 2020 3360
rect 2070 3352 2112 3360
rect 2070 3328 2078 3352
rect 2102 3328 2112 3352
rect 2070 3320 2112 3328
rect 2289 3332 2332 3340
rect 1990 3274 2032 3280
rect 1990 3251 1999 3274
rect 2021 3251 2032 3274
rect 1990 3242 2032 3251
rect 1945 3212 1986 3221
rect 2081 3220 2110 3320
rect 2289 3300 2298 3332
rect 2324 3300 2332 3332
rect 2289 3290 2332 3300
rect 1945 3030 1952 3212
rect 1978 3030 1986 3212
rect 1945 2996 1986 3030
rect 2070 3211 2110 3220
rect 2070 3029 2077 3211
rect 2103 3029 2110 3211
rect 2070 2996 2110 3029
<< via1 >>
rect 1766 3954 1793 3987
rect 1627 3827 1653 3853
rect 1887 3797 1913 3823
rect 1766 3652 1793 3685
rect 2076 3650 2103 3987
rect 2281 4005 2316 4031
rect 2467 3996 2493 4022
rect 1592 3372 1618 3399
rect 1766 3370 1792 3396
rect 2366 3430 2392 3456
rect 2298 3388 2324 3414
rect 1888 3298 1914 3324
rect 2298 3300 2324 3332
rect 1952 3030 1978 3212
<< metal2 >>
rect 2256 4031 2340 4038
rect 1760 3987 1800 4013
rect 1760 3954 1766 3987
rect 1793 3954 1800 3987
rect 1760 3929 1800 3954
rect 2070 3987 2110 4025
rect 2256 4005 2281 4031
rect 2316 4005 2340 4031
rect 2256 3998 2340 4005
rect 2460 4022 2500 4030
rect 1760 3860 1790 3929
rect 2070 3860 2076 3987
rect 1620 3853 2076 3860
rect 1620 3827 1627 3853
rect 1653 3827 2076 3853
rect 1620 3820 1660 3827
rect 1760 3711 1790 3827
rect 1879 3823 1921 3827
rect 1879 3797 1887 3823
rect 1913 3797 1921 3823
rect 1879 3789 1921 3797
rect 1760 3685 1800 3711
rect 1760 3652 1766 3685
rect 1793 3652 1800 3685
rect 1760 3627 1800 3652
rect 2070 3650 2076 3827
rect 2103 3860 2110 3987
rect 2290 3860 2320 3998
rect 2460 3996 2467 4022
rect 2493 3996 2500 4022
rect 2460 3990 2500 3996
rect 2103 3827 2320 3860
rect 2103 3650 2110 3827
rect 2070 3625 2110 3650
rect 2290 3422 2320 3827
rect 2356 3456 2400 3466
rect 2356 3430 2366 3456
rect 2392 3450 2400 3456
rect 2470 3450 2500 3990
rect 2392 3430 2500 3450
rect 2289 3414 2333 3422
rect 2356 3420 2500 3430
rect 1580 3400 1630 3410
rect 1759 3400 1800 3405
rect 1580 3399 1800 3400
rect 1580 3372 1592 3399
rect 1618 3396 1800 3399
rect 1618 3372 1766 3396
rect 1580 3370 1766 3372
rect 1792 3370 1800 3396
rect 2289 3388 2298 3414
rect 2324 3388 2333 3414
rect 2289 3380 2333 3388
rect 1580 3360 1630 3370
rect 1680 3320 1710 3370
rect 1759 3362 1800 3370
rect 2289 3332 2332 3340
rect 1880 3324 1922 3332
rect 1880 3320 1888 3324
rect 1680 3298 1888 3320
rect 1914 3320 1922 3324
rect 2289 3320 2298 3332
rect 1914 3300 2298 3320
rect 2324 3300 2332 3332
rect 1914 3298 2332 3300
rect 1680 3290 2332 3298
rect 1945 3221 1975 3290
rect 1945 3212 1986 3221
rect 1945 3030 1952 3212
rect 1978 3030 1986 3212
rect 1945 2996 1986 3030
<< labels >>
rlabel locali 2378 3186 2410 3200 1 cp
rlabel metal1 1637 3487 1691 3502 1 dn
rlabel locali 1871 4378 1899 4393 1 gnd!
rlabel metal1 1683 4140 1711 4155 1 up
rlabel locali 1659 3778 1687 3793 1 vdd
<< end >>
