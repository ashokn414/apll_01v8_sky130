***inverter circuit***
.param L=0.15
.param W=0.42
.include "sky130_fd_pr/models/corners/tt.spice"

X1 out in GND GND sky130_fd_pr__nfet_01v8 l={L} w={W}
X2 VDD in out VDD sky130_fd_pr__pfet_01v8 l={L} w={2.5*W}

***set gnd and power***
 
Vdd VDD 0 1.8
Vin in 0 0 pulse(0 1.8 0 10p 10p 1n 2n) 

.op
.tran 10p 4n
.end

