***charge_pump circuit***
.param L=0.15
.param W=0.42
.include "/home/ashok/sky130_fd_pr/models/corners/tt.spice"

***netlist for charge pump***
X7 UP_bar UP 0 0 sky130_fd_pr__nfet_01v8 l={L} w={W}
X8 DOWN_bar Down 0 0 sky130_fd_pr__nfet_01v8 l={L} w={W}
X12 VDD Down DOWN_bar VDD sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X14 VDD UP UP_bar VDD sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X15 UP_bar 0 N001 N001 sky130_fd_pr__nfet_01v8 l={L} w={W}
X16 DOWN_bar 0 N004 N004 sky130_fd_pr__nfet_01v8 l={L} w={W}
X17 N003 N004 N003 N003 sky130_fd_pr__nfet_01v8 l={L} w={W}
X18 0 VDD VDD 0 sky130_fd_pr__nfet_01v8 l={L} w={W}
X19 CP VDD N003 N003 sky130_fd_pr__nfet_01v8 l={L} w={W}
X20 N003 Down 0 0 sky130_fd_pr__nfet_01v8 l={L} w={55*W}
X21 N001 VDD UP_bar N001 sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X22 N004 VDD DOWN_bar N004 sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X23 N002 UP N002 N002 sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X24 0 0 VDD VDD sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X25 N002 0 CP N002 sky130_fd_pr__pfet_01v8 l={L} w={3*W}
X26 VDD N001 N002 VDD sky130_fd_pr__pfet_01v8 l={L} w={166*W}
V1 VDD 0 1.8

***set power***
up1 UP 0 0 pulse(0 1.8 0 10p 10p 1n 5n)
do1 Down 0 0 pulse(0 1.8 0 10p 10p 1n 7n)

.op
.tran 10p 50n
.end
