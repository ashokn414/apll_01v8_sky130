inverter circuit
.param L=0.15
.param W=0.42
.include "/home/ashok/sky130_fd_pr/models/corners/tt.spice"
* instantiate the inverter
Xinv Y A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_1
* SPICE3 file created from sky130_fd_sc_hd__inv_1.ext - technology:sky130A
.subckt sky130_fd_sc_hd__inv_1 Y A VPB VNB VGND VPWR
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 w={2*W} l={L}
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w={2*W} l={L}
.ends
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8
* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 2n
.control
run
plot A Y i(Vin)
.endc
.end
