***inv_20_10 circuit***
.param L=0.15
.param W=0.42
.include "/home/ashok/sky130_fd_pr/models/corners/tt.spice"

X1 Out In 0 0 sky130_fd_pr__nfet_01v8 l={L} w={2*W}
X2 Out In N001 N001 sky130_fd_pr__pfet_01v8 l={L} w={4*W}
V1 N001 0 1.8
***set gnd and power***
 
Vin In 0 0 pulse(0 1.8 0 10p 10p 1n 2n) 

.op
.tran 10p 4n
.end

