* /home/shabari/esim/esim-1.1.3/src/subcircuitlibrary/testinv/testinv.cir
.param L=0.15
.param W=0.42
.include "sky130_fd_pr/models/corners/tt.spice"
X1 N001 B 0 0 sky130_fd_pr__nfet_01v8 l=L w=W
X2 NAND A N001 NC_01 sky130_fd_pr__nfet_01v8 l=L w=W
X3 AND Abar 0 0 sky130_fd_pr__nfet_01v8 l=L w=W
X4 AND Bbar 0 0 sky130_fd_pr__nfet_01v8 l=L w=W
X5 VDD AND NAND VDD sky130_fd_pr__pfet_01v8 l=L w=W
X6 VDD NAND AND VDD sky130_fd_pr__pfet_01v8 l=L w=W
X7 VDD B Bbar VDD sky130_fd_pr__pfet_01v8 l=L w=W
X8 VDD A Abar VDD sky130_fd_pr__pfet_01v8 l=L w=W
X9 Abar A 0 0 sky130_fd_pr__nfet_01v8 l=L w=W
X10 Bbar B 0 0 sky130_fd_pr__nfet_01v8 l=L w=W
V1 VDD 0 2.5
V2 A 0 PULSE(0 2.5 0 100ps 100ps 20n 40n)
V3 B 0 PULSE(0 2.5 0 100ps 100ps 40n 80n)

.tran 10p 80n

.end



