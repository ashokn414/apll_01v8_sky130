* NGSPICE file created from vco.ext - technology: sky130A


* Top level circuit vco

X0 a_915_n134# a_100_n200# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X1 a_540_n411# a_330_n411# a_495_n411# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_705_n411# vin gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_495_n411# vin gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_100_n200# a_100_n200# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X5 a_330_n411# a_280_n277# a_285_n411# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_285_n411# vin gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_960_n411# a_750_n411# a_915_n134# vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X8 a_705_n134# a_100_n200# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X9 a_750_n411# a_540_n411# a_705_n134# vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 vout a_280_n277# gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_540_n411# a_330_n411# a_495_n134# vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 a_1125_n411# vin gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_495_n134# a_100_n200# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X14 a_330_n411# a_280_n277# a_285_n134# vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_285_n134# a_100_n200# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X16 a_280_n277# a_960_n411# a_1125_n411# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 vout a_280_n277# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X18 a_1125_n134# a_100_n200# vdd vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X19 a_915_n411# vin gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_100_n200# vin gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_280_n277# a_960_n411# a_1125_n134# vdd sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X22 a_960_n411# a_750_n411# a_915_n411# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_750_n411# a_540_n411# a_705_n411# gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.end

